    (** * Examples of Stable Category Theory Structures

        This module provides concrete trivial and non-trivial examples for the abstract structures
        defined in our formalization, built incrementally from the simplest
        to more complex. The purpose of the trivial examples is to establish non-vacuity.
    *)

    From HoTT Require Import Basics Types Categories.
    From HoTT.Categories Require Import Category.

    Require Import ZeroObjects.

    (** * Example 1: The Simplest Zero Object *)

    Module SimplestZeroObject.

      (** The one-object, one-morphism category. *)
      Definition OneCat : PreCategory.
      Proof.
        simple refine (@Build_PreCategory
          Unit                          (* Type of objects *)
          (fun _ _ => Unit)            (* Morphism type *)
          (fun _ => tt)                (* Identity *)
          (fun _ _ _ _ _ => tt)        (* Composition *)
          _ _ _ _).                    
        - (* associativity *)
          intros s d d' d'' m1 m2 m3.
          destruct m1, m2, m3.
          reflexivity.
        - (* left identity *)  
          intros a b f.
          destruct a, b, f.
          reflexivity.
        - (* right identity *)
          intros a b f.
          destruct a, b, f.
          reflexivity.
      Defined.

        (** The unique object is a zero object. *)
        Theorem one_object_is_zero : ZeroObject OneCat.
        Proof.
          simple refine (Build_ZeroObject OneCat tt _ _).
        Defined.

      (** Verify the zero morphism is what we expect. *)
      Lemma zero_morphism_is_tt : 
        zero_morphism one_object_is_zero tt tt = tt.
      Proof.
        reflexivity.
      Qed.

    End SimplestZeroObject.

    (** * Example 2: A Category with Biproducts *)

    Module SimpleBiproductCategory.

    Require Import Biproducts.

      (** A two-object category with biproducts. 
          Objects: {0, 1} where 0 is zero object
          Morphisms: only identities and unique morphisms to/from 0 *)
      
      Inductive TwoObj : Type := Zero | One.
      
      Definition TwoMor (X Y : TwoObj) : Type :=
        match X, Y with
        | Zero, _ => Unit    (* unique morphism from zero *)
        | _, Zero => Unit    (* unique morphism to zero *)
        | One, One => Unit   (* identity on One *)
        end.
      
      Definition two_id (X : TwoObj) : TwoMor X X :=
        match X with
        | Zero => tt
        | One => tt
        end.
      
      Definition two_comp {X Y Z : TwoObj} (g : TwoMor Y Z) (f : TwoMor X Y) : TwoMor X Z.
      Proof.
        destruct X, Y, Z; try exact tt.
      Defined.
      
    Definition TwoCat : PreCategory.
    Proof.
      simple refine (@Build_PreCategory
        TwoObj
        TwoMor
        two_id
        (@two_comp)
        _ _ _ _).
      - (* associativity *)
        intros s d d' d'' m1 m2 m3.
        destruct s, d, d', d''; 
        try destruct m1; try destruct m2; try destruct m3; 
        reflexivity.
      - (* left identity *)
        intros a b f.
        destruct a, b; destruct f; reflexivity.
      - (* right identity *)
        intros a b f.
        destruct a, b; destruct f; reflexivity.
      - (* truncation: morphisms form a set *)
        intros s d.
        destruct s, d; apply _.
    Defined.
      
    (** Zero is the zero object. *)
    Theorem two_zero : ZeroObject TwoCat.
    Proof.
      simple refine (Build_ZeroObject TwoCat Zero _ _).
      - (* Zero is initial: unique morphism from Zero to any Y *)
        intro Y.
        destruct Y.
        + (* Y = Zero *)
          apply Build_Contr with (center := tt).
          intro f.
          unfold morphism in f; simpl in f.
          destruct f; reflexivity.
        + (* Y = One *)
          apply Build_Contr with (center := tt).
          intro f.
          unfold morphism in f; simpl in f.
          destruct f; reflexivity.
    Defined.
      
    (** The biproduct of One and One exists (it's One). *)
    Definition one_plus_one : @Biproduct TwoCat One One two_zero.
    Proof.
      (* Biproduct data *)
      pose (bdata := Build_BiproductData TwoCat One One One tt tt tt tt).
      
      (* Biproduct axioms *)
      assert (bis : IsBiproduct bdata two_zero).
      {
        simple refine (Build_IsBiproduct _ _ _ _ _ _ _ _ _).
        - reflexivity.  (* outl ∘ inl = id *)
        - reflexivity.  (* outr ∘ inr = id *)
        - reflexivity.  (* outl ∘ inr = 0 *)
        - reflexivity.  (* outr ∘ inl = 0 *)
      }
      

    (* Universal property *)
    assert (buni : HasBiproductUniversal bdata).
    {
      simple refine (Build_HasBiproductUniversal _ _ _ _ _ _).
      - (* Coproduct universal *)
        intros Z f g.
        destruct Z.
        + (* Z = Zero *)
          destruct f, g.
          apply Build_Contr with (center := (tt; (idpath, idpath))).
          intros [h' [p q]].
          apply path_sigma_uncurried.
          exists (match h' with tt => idpath end).
          simpl.
          apply path_prod; apply path_ishprop.
        + (* Z = One *)
          destruct f, g.
          apply Build_Contr with (center := (tt; (idpath, idpath))).
          intros [h' [p q]].
          apply path_sigma_uncurried.
          exists (match h' with tt => idpath end).
          simpl.
          apply path_prod; apply path_ishprop.
      - (* Product universal *)
        intros Z f g.
        destruct Z.
        + (* Z = Zero *)
          destruct f, g.
          apply Build_Contr with (center := (tt; (idpath, idpath))).
          intros [h' [p q]].
          apply path_sigma_uncurried.
          exists (match h' with tt => idpath end).
          simpl.
          apply path_prod; apply path_ishprop.
        + (* Z = One *)
          destruct f, g.
          apply Build_Contr with (center := (tt; (idpath, idpath))).
          intros [h' [p q]].
          apply path_sigma_uncurried.
          exists (match h' with tt => idpath end).
          simpl.
          apply path_prod; apply path_ishprop.
    }
  exact (Build_Biproduct _ _ _ _ bdata bis buni).
    Defined.

  End SimpleBiproductCategory.

  Module TwoCatAdditive.
    Import SimpleBiproductCategory.
    Require Import Biproducts.
    Require Import AdditiveCategories.
    
    (* First prove all biproducts exist *)
    Definition two_all_biproducts (X Y : object TwoCat) : Biproduct X Y two_zero.
    Proof.
      destruct X, Y.
      - (* Zero ⊕ Zero = Zero *)
        pose (bdata := Build_BiproductData TwoCat Zero Zero Zero tt tt tt tt).
  assert (bis : IsBiproduct bdata two_zero).
        {
          simple refine (Build_IsBiproduct _ _ _ _ _ _ _ _ _).
          - (* outl ∘ inl = id *) reflexivity.
          - (* outr ∘ inr = id *) reflexivity.
          - (* outl ∘ inr = 0 *) reflexivity.
          - (* outr ∘ inl = 0 *) reflexivity.
        }
  assert (buni : HasBiproductUniversal bdata).
        {
          simple refine (Build_HasBiproductUniversal _ _ _ _ _ _).
          - (* Coproduct universal *)
            intros W f g.
            destruct W.
            + (* W = Zero *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
            + (* W = One *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
  }
        exact (Build_Biproduct _ _ _ _ bdata bis buni).
  - (* Zero ⊕ One = One *)
        pose (bdata := Build_BiproductData TwoCat Zero One One tt tt tt tt).
        assert (bis : IsBiproduct bdata two_zero).
        {
          simple refine (Build_IsBiproduct _ _ _ _ _ _ _ _ _).
          - (* outl ∘ inl = id *) reflexivity.
          - (* outr ∘ inr = id *) reflexivity.
          - (* outl ∘ inr = 0 *) reflexivity.
          - (* outr ∘ inl = 0 *) reflexivity.
        }
  assert (buni : HasBiproductUniversal bdata).
        {
          simple refine (Build_HasBiproductUniversal _ _ _ _ _ _).
          - (* Coproduct universal *)
            intros W f g.
            destruct W.
            + (* W = Zero *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
            + (* W = One *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
  - (* Product universal *)
            intros W f g.
            destruct W.
            + (* W = Zero *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
            + (* W = One *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
        }
        exact (Build_Biproduct _ _ _ _ bdata bis buni).
  - (* One ⊕ Zero = One *)
        pose (bdata := Build_BiproductData TwoCat One Zero One tt tt tt tt).
        assert (bis : IsBiproduct bdata two_zero).
        {
          simple refine (Build_IsBiproduct _ _ _ _ _ _ _ _ _).
          - (* outl ∘ inl = id *) reflexivity.
          - (* outr ∘ inr = id *) reflexivity.
          - (* outl ∘ inr = 0 *) reflexivity.
          - (* outr ∘ inl = 0 *) reflexivity.
        }
  assert (buni : HasBiproductUniversal bdata).
        {
          simple refine (Build_HasBiproductUniversal _ _ _ _ _ _).
          - (* Coproduct universal *)
            intros W f g.
            destruct W.
            + (* W = Zero *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
            + (* W = One *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
          - (* Product universal *)
            intros W f g.
            destruct W.
            + (* W = Zero *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
            + (* W = One *)
              destruct f, g.
              apply Build_Contr with (center := (tt; (idpath, idpath))).
              intros [h' [p q]].
              apply path_sigma_uncurried.
              exists (match h' with tt => idpath end).
              simpl.
              apply path_prod; apply path_ishprop.
        }
        exact (Build_Biproduct _ _ _ _ bdata bis buni).
  - (* One ⊕ One = One *)
        exact one_plus_one.
    Defined.

  Definition TwoAdditive : AdditiveCategory.
    Proof.
      exact (Build_AdditiveCategory TwoCat two_zero two_all_biproducts).
    Defined.

  End TwoCatAdditive.

  Module ChainComplexExample.
    From HoTT Require Import Basics Types.
    Require Import ZeroObjects Biproducts AdditiveCategories PreStableCategories.
    
    Section ChainComplexes.
      Context `{Funext}.
      
      (* First, we need abelian groups *)
      Record AbelianGroup : Type := {
        carrier : Type;
        zero : carrier;
        plus : carrier -> carrier -> carrier;
        neg : carrier -> carrier
      }.
      
      (* Group axioms *)
      Record AbelianGroup_laws (G : AbelianGroup) : Type := {
        plus_assoc : forall x y z : carrier G, 
          plus G x (plus G y z) = plus G (plus G x y) z;
        plus_zero_l : forall x : carrier G, plus G (zero G) x = x;
        plus_zero_r : forall x : carrier G, plus G x (zero G) = x;
        plus_neg_l : forall x : carrier G, plus G (neg G x) x = zero G;
        plus_neg_r : forall x : carrier G, plus G x (neg G x) = zero G;
        plus_comm : forall x y : carrier G, plus G x y = plus G y x
      }.
      
      (* Complete abelian group with laws and set requirement *)
      Record AbelianGroupWithLaws : Type := {
        group : AbelianGroup;
        laws : AbelianGroup_laws group;
        carrier_is_set : IsHSet (carrier group)
      }.
      
      (* Group homomorphisms *)
      Record GroupHom (G H : AbelianGroupWithLaws) : Type := {
        hom_map : carrier (group G) -> carrier (group H);
        hom_zero : hom_map (zero (group G)) = zero (group H);
        hom_plus : forall x y : carrier (group G), 
          hom_map (plus (group G) x y) = plus (group H) (hom_map x) (hom_map y)
      }.
      
      (* Helper: In a set, all paths between two elements are equal *)
      Lemma path_hset {A : Type} {HSet : IsHSet A} (x y : A) (p q : x = y) : p = q.
      Proof.
        apply path_ishprop.
      Qed.

    (* Identity homomorphism *)
      Definition id_hom (G : AbelianGroupWithLaws) : GroupHom G G.
      Proof.
        refine (Build_GroupHom G G (fun x => x) _ _).
        - (* hom_zero *) reflexivity.
        - (* hom_plus *) intros x y. reflexivity.
      Defined.

  (* Helper: In an HSet, all paths between two elements are equal *)
      Lemma hset_path_unique {A : Type} (HA : IsHSet A) {x y : A} (p q : x = y) : p = q.
      Proof.
        apply path_ishprop.
      Qed.

  (* Two homomorphisms are equal if their underlying functions are equal *)
      Lemma GroupHom_eq {G K : AbelianGroupWithLaws} (f g : GroupHom G K) :
        hom_map G K f = hom_map G K g -> f = g.
      Proof.
        intro p.
        destruct f as [f_map f_zero f_plus].
        destruct g as [g_map g_zero g_plus].
        simpl in p.
        destruct p.
        (* Now f_map = g_map definitionally *)
        assert (Hz : f_zero = g_zero).
        {
          apply hset_path_unique.
          apply (carrier_is_set K).
        }
        assert (Hp : f_plus = g_plus).
        {
          apply path_forall; intro x.
          apply path_forall; intro y.
          apply hset_path_unique.
          apply (carrier_is_set K).
        }
        destruct Hz, Hp.
        reflexivity.
      Qed.

  (* Composition of homomorphisms *)
      Definition comp_hom {A B C : AbelianGroupWithLaws} 
        (g : GroupHom B C) (f : GroupHom A B) : GroupHom A C.
      Proof.
        refine (Build_GroupHom A C 
          (fun x => hom_map B C g (hom_map A B f x)) _ _).
        - (* hom_zero *)
          rewrite (hom_zero A B f).
          rewrite (hom_zero B C g).
          reflexivity.
        - (* hom_plus *)
          intros x y.
          rewrite (hom_plus A B f).
          rewrite (hom_plus B C g).
          reflexivity.
      Defined.

  (* The property of being a group homomorphism is a proposition *)
      Lemma IsGroupHom_HProp (A B : AbelianGroupWithLaws) 
        (f : carrier (group A) -> carrier (group B)) :
        IsHProp ((f (zero (group A)) = zero (group B)) * 
                 (forall x y, f (plus (group A) x y) = plus (group B) (f x) (f y))).
      Proof.
        (* First show the components are props *)
        assert (H1 : IsHProp (f (zero (group A)) = zero (group B))).
        { 
          apply hprop_allpath.
          intros p q.
          apply hset_path_unique.
          apply (carrier_is_set B).
        }
        assert (H2 : IsHProp (forall x y, f (plus (group A) x y) = plus (group B) (f x) (f y))).
        {
          apply hprop_allpath.
          intros p q.
          apply path_forall. intro x.
          apply path_forall. intro y.
          apply hset_path_unique.
          apply (carrier_is_set B).
        }
        (* Now the product *)
        apply istrunc_prod; assumption.
      Qed.

  (* GroupHom is equivalent to a sigma type *)
      Definition GroupHom_to_sig (A B : AbelianGroupWithLaws) (h : GroupHom A B) :
        {f : carrier (group A) -> carrier (group B) & 
         (f (zero (group A)) = zero (group B)) * 
         (forall x y, f (plus (group A) x y) = plus (group B) (f x) (f y))}.
      Proof.
        exists (hom_map A B h).
        split.
        - apply (hom_zero A B h).
        - apply (hom_plus A B h).
      Defined.

  (* Sigma type to GroupHom *)
      Definition sig_to_GroupHom (A B : AbelianGroupWithLaws) 
        (s : {f : carrier (group A) -> carrier (group B) & 
              (f (zero (group A)) = zero (group B)) * 
              (forall x y, f (plus (group A) x y) = plus (group B) (f x) (f y))}) 
        : GroupHom A B.
      Proof.
        destruct s as [f [hz hp]].
        exact (Build_GroupHom A B f hz hp).
      Defined.

  (* They are inverses *)
      Lemma GroupHom_sig_equiv_sect (A B : AbelianGroupWithLaws) (h : GroupHom A B) :
        sig_to_GroupHom A B (GroupHom_to_sig A B h) = h.
      Proof.
        destruct h as [f hz hp].
        reflexivity.
      Qed.

  (* The other inverse *)
      Lemma GroupHom_sig_equiv_retr (A B : AbelianGroupWithLaws) 
        (s : {f : carrier (group A) -> carrier (group B) & 
              (f (zero (group A)) = zero (group B)) * 
              (forall x y, f (plus (group A) x y) = plus (group B) (f x) (f y))}) :
        GroupHom_to_sig A B (sig_to_GroupHom A B s) = s.
      Proof.
        destruct s as [f [hz hp]].
        reflexivity.
      Qed.

  (* The equivalence *)
      Definition GroupHom_sig_equiv (A B : AbelianGroupWithLaws) :
        GroupHom A B <~> 
        {f : carrier (group A) -> carrier (group B) & 
         (f (zero (group A)) = zero (group B)) * 
         (forall x y, f (plus (group A) x y) = plus (group B) (f x) (f y))}.
      Proof.
        apply (equiv_adjointify 
          (GroupHom_to_sig A B)
          (sig_to_GroupHom A B)).
        - intro s. apply GroupHom_sig_equiv_retr.
        - intro h. apply GroupHom_sig_equiv_sect.
      Defined.

  (* Helper: Function types are HSets when codomain is *)
  Lemma fun_is_hset `{Funext} (A B : Type) (HB : IsHSet B) : IsHSet (A -> B).
  Proof.
    change (IsTrunc 0 (A -> B)).
    apply istrunc_forall.
  Qed.

  (* Helper: Product types are HSets when both components are *)
  Lemma prod_is_hset (A B : Type) (HA : IsHSet A) (HB : IsHSet B) : IsHSet (A * B).
  Proof.
    apply istrunc_prod; assumption.
  Qed.

  (* Helper: Sigma types are HSets when base is HSet and fibers are HProps *)
  Lemma sig_is_hset_from_hprop (A : Type) (P : A -> Type) 
    (HA : IsHSet A) (HP : forall a, IsHProp (P a)) : IsHSet (sig P).
  Proof.
    apply istrunc_sigma.
  Qed.

  (* Helper: Paths in sets are HProps *)
  Lemma path_ishprop_hset (A : Type) (HA : IsHSet A) (x y : A) : IsHProp (x = y).
  Proof.
    exact (HA x y).
  Qed.

  (* Helper: Product of HProps is HProp *)
  Lemma prod_hprop (A B : Type) (HA : IsHProp A) (HB : IsHProp B) : IsHProp (A * B).
  Proof.
    change (IsTrunc (-1) (A * B)).
    apply istrunc_prod; assumption.
  Qed.

  (* Helper: Forall over HProps is HProp *)
  Lemma forall_hprop `{Funext} (A : Type) (P : A -> Type) 
    (HP : forall a, IsHProp (P a)) : IsHProp (forall a, P a).
  Proof.
    change (IsTrunc (-1) (forall a, P a)).
    apply istrunc_forall.
  Qed.

  (* Helper: The GroupHom property is an HProp for any function *)
  Lemma GroupHom_property_is_hprop `{Funext} (A B : AbelianGroupWithLaws) 
    (f : carrier (group A) -> carrier (group B)) :
    IsHProp ((f (zero (group A)) = zero (group B)) * 
             (forall x y, f (plus (group A) x y) = plus (group B) (f x) (f y))).
  Proof.
    apply prod_hprop.
    - (* First component is HProp *)
      apply path_ishprop_hset.
      apply (carrier_is_set B).
    - (* Second component is HProp *)
      apply forall_hprop. intro x.
      apply forall_hprop. intro y.
      apply path_ishprop_hset.
      apply (carrier_is_set B).
  Qed.

  (* Now we can prove GroupHom is an HSet *)
  Global Instance GroupHom_IsHSet `{Funext} (A B : AbelianGroupWithLaws) : IsHSet (GroupHom A B).
  Proof.
    (* First show the sigma type is an HSet *)
    assert (HSig : IsHSet {f : carrier (group A) -> carrier (group B) & 
                           (f (zero (group A)) = zero (group B)) * 
                           (forall x y, f (plus (group A) x y) = plus (group B) (f x) (f y))}).
    {
      apply sig_is_hset_from_hprop.
      - (* Base type is HSet *)
        apply fun_is_hset.
        apply (carrier_is_set B).
      - (* Fibers are HProps *)
        intro f.
        apply GroupHom_property_is_hprop.
    }
    (* Now use the equivalence *)
    exact (istrunc_equiv_istrunc _ (GroupHom_sig_equiv A B)^-1).
  Qed.

  (* The zero homomorphism *)
  Definition zero_hom (A B : AbelianGroupWithLaws) : GroupHom A B.
  Proof.
    refine (Build_GroupHom A B (fun _ => zero (group B)) _ _).
    - (* hom_zero *) reflexivity.
    - (* hom_plus *) 
      intros x y.
      symmetry.
      apply (plus_zero_l (group B) (laws B)).
  Defined.

  (* Composition is associative *)
  Lemma comp_hom_assoc {A B C D : AbelianGroupWithLaws}
    (h : GroupHom C D) (g : GroupHom B C) (f : GroupHom A B) :
    comp_hom h (comp_hom g f) = comp_hom (comp_hom h g) f.
  Proof.
    apply GroupHom_eq.
    reflexivity.
  Qed.

  (* Composition with identity on the left *)
  Lemma comp_hom_id_left {A B : AbelianGroupWithLaws} (f : GroupHom A B) :
    comp_hom (id_hom B) f = f.
  Proof.
    apply GroupHom_eq.
    reflexivity.
  Qed.

  (* Composition with identity on the right *)
  Lemma comp_hom_id_right {A B : AbelianGroupWithLaws} (f : GroupHom A B) :
    comp_hom f (id_hom A) = f.
  Proof.
    apply GroupHom_eq.
    reflexivity.
  Qed.

  (* The category of abelian groups *)
  Definition AbGroupCat `{Funext} : PreCategory.
  Proof.
    refine (@Build_PreCategory
      AbelianGroupWithLaws
      GroupHom
      id_hom
      (fun A B C => comp_hom)
      _ _ _ _).
    - (* associativity *)
      intros A B C D f g h.
      symmetry.
      apply comp_hom_assoc.
    - (* left identity *)
      intros A B f.
      apply comp_hom_id_left.
    - (* right identity *)
      intros A B f.
      apply comp_hom_id_right.
  Defined.

  (* The trivial abelian group *)
  Definition TrivialGroup : AbelianGroupWithLaws.
  Proof.
    refine (Build_AbelianGroupWithLaws
      (Build_AbelianGroup Unit tt (fun _ _ => tt) (fun _ => tt))
      _ _).
    - (* laws *)
      refine (Build_AbelianGroup_laws _ _ _ _ _ _ _).
      + (* plus_assoc *) intros x y z. destruct x, y, z. reflexivity.
      + (* plus_zero_l *) intros x. destruct x. reflexivity.
      + (* plus_zero_r *) intros x. destruct x. reflexivity.
      + (* plus_neg_l *) intros x. destruct x. reflexivity.
      + (* plus_neg_r *) intros x. destruct x. reflexivity.
      + (* plus_comm *) intros x y. destruct x, y. reflexivity.
  Defined.

  (* TrivialGroup is the zero object in AbGroupCat *)
  Theorem TrivialGroup_is_zero : ZeroObject AbGroupCat.
  Proof.
    refine (Build_ZeroObject AbGroupCat TrivialGroup _ _).
    - (* initial *)
      intro X.
      simple refine (Build_Contr _ _ _).
      + (* center: the zero morphism *)
        simple refine (Build_GroupHom TrivialGroup X (fun _ => zero (group X)) _ _).
        * (* hom_zero *)
          reflexivity.
        * (* hom_plus *)
          intros x y.
          simpl.
          symmetry.
          apply (plus_zero_l (group X) (laws X)).
      + (* contr: uniqueness *)
        intro f.
        apply GroupHom_eq.
        apply path_forall. intro x.
        destruct x.
        simpl.
        symmetry.
        exact (hom_zero TrivialGroup X f).
    - (* terminal *)
      intro X.
      simple refine (Build_Contr _ _ _).
      + (* center *)
        simple refine (Build_GroupHom X TrivialGroup (fun _ => tt) _ _).
        * (* hom_zero *)
          reflexivity.
        * (* hom_plus *)
          intros x y. reflexivity.
      + (* contr: uniqueness *)
        intro f.
        apply GroupHom_eq.
        apply path_forall. intro x.
        destruct (hom_map X TrivialGroup f x).
        reflexivity.
  Defined.

  (* Direct sum of abelian groups *)
  Definition DirectSum (A B : AbelianGroupWithLaws) : AbelianGroupWithLaws.
  Proof.
    refine (Build_AbelianGroupWithLaws
      (Build_AbelianGroup 
        (carrier (group A) * carrier (group B))
        (zero (group A), zero (group B))
        (fun p1 p2 => (plus (group A) (fst p1) (fst p2), 
                       plus (group B) (snd p1) (snd p2)))
        (fun p => (neg (group A) (fst p), neg (group B) (snd p))))
      _ _).
    - (* laws *)
      refine (Build_AbelianGroup_laws _ _ _ _ _ _ _).
      + (* plus_assoc *)
        intros [a1 b1] [a2 b2] [a3 b3].
        simpl.
        f_ap.
        * apply (plus_assoc (group A) (laws A)).
        * apply (plus_assoc (group B) (laws B)).
      + (* plus_zero_l *)
        intros [a b].
        simpl.
        f_ap.
        * apply (plus_zero_l (group A) (laws A)).
        * apply (plus_zero_l (group B) (laws B)).
      + (* plus_zero_r *)
        intros [a b].
        simpl.
        f_ap.
        * apply (plus_zero_r (group A) (laws A)).
        * apply (plus_zero_r (group B) (laws B)).
      + (* plus_neg_l *)
        intros [a b].
        simpl.
        f_ap.
        * apply (plus_neg_l (group A) (laws A)).
        * apply (plus_neg_l (group B) (laws B)).
      + (* plus_neg_r *)
        intros [a b].
        simpl.
        f_ap.
        * apply (plus_neg_r (group A) (laws A)).
        * apply (plus_neg_r (group B) (laws B)).
      + (* plus_comm *)
        intros [a1 b1] [a2 b2].
        simpl.
        f_ap.
        * apply (plus_comm (group A) (laws A)).
        * apply (plus_comm (group B) (laws B)).
    - (* carrier_is_set *)
      apply prod_is_hset.
      + apply (carrier_is_set A).
      + apply (carrier_is_set B).
  Defined.

  (* First projection from direct sum *)
  Definition proj1 (A B : AbelianGroupWithLaws) : GroupHom (DirectSum A B) A.
  Proof.
    refine (Build_GroupHom (DirectSum A B) A fst _ _).
    - (* hom_zero *)
      reflexivity.
    - (* hom_plus *)
      intros [a1 b1] [a2 b2].
      reflexivity.
  Defined.

  (* Second projection from direct sum *)
  Definition proj2 (A B : AbelianGroupWithLaws) : GroupHom (DirectSum A B) B.
  Proof.
    refine (Build_GroupHom (DirectSum A B) B snd _ _).
    - (* hom_zero *)
      reflexivity.
    - (* hom_plus *)
      intros [a1 b1] [a2 b2].
      reflexivity.
  Defined.

  (* First injection into direct sum *)
  Definition inj1 (A B : AbelianGroupWithLaws) : GroupHom A (DirectSum A B).
  Proof.
    refine (Build_GroupHom A (DirectSum A B) (fun a => (a, zero (group B))) _ _).
    - (* hom_zero *)
      reflexivity.
    - (* hom_plus *)
      intros a1 a2.
      simpl.
      f_ap.
      symmetry.
      apply (plus_zero_l (group B) (laws B)).
  Defined.

  (* Second injection into direct sum *)
  Definition inj2 (A B : AbelianGroupWithLaws) : GroupHom B (DirectSum A B).
  Proof.
    refine (Build_GroupHom B (DirectSum A B) (fun b => (zero (group A), b)) _ _).
    - (* hom_zero *)
      reflexivity.
    - (* hom_plus *)
      intros b1 b2.
      simpl.
      f_ap.
      symmetry.
      apply (plus_zero_l (group A) (laws A)).
  Defined.

  (* Chain complexes over abelian groups *)
  Record ChainComplex := {
    ob : nat -> AbelianGroupWithLaws;
    diff : forall n, GroupHom (ob (S n)) (ob n);
    diff_squared : forall n, 
      comp_hom (diff n) (diff (S n)) = zero_hom (ob (S (S n))) (ob n)
  }.

  (* Chain maps between chain complexes *)
  Record ChainMap (C D : ChainComplex) := {
    map_ob : forall n, GroupHom (ob C n) (ob D n);
    map_commutes : forall n,
      comp_hom (map_ob n) (diff C n) = comp_hom (diff D n) (map_ob (S n))
  }.

  (* Identity chain map *)
  Definition id_chain_map (C : ChainComplex) : ChainMap C C.
  Proof.
    refine (Build_ChainMap C C (fun n => id_hom (ob C n)) _).
    intro n.
    rewrite comp_hom_id_left.
    rewrite comp_hom_id_right.
    reflexivity.
  Defined.

   (* Composition of chain maps *)
  Definition comp_chain_map {A B C : ChainComplex} 
    (g : ChainMap B C) (f : ChainMap A B) : ChainMap A C.
  Proof.
    refine (Build_ChainMap A C 
      (fun n => comp_hom (map_ob B C g n) (map_ob A B f n)) _).
    intro n.
    rewrite <- comp_hom_assoc.
    rewrite (map_commutes A B f n).
    rewrite comp_hom_assoc.
    rewrite (map_commutes B C g n).
    rewrite <- comp_hom_assoc.
    reflexivity.
  Defined.

  (* Chain maps are equal if their components are equal *)
  Lemma ChainMap_eq {C D : ChainComplex} (f g : ChainMap C D) :
    (forall n, map_ob C D f n = map_ob C D g n) -> f = g.
  Proof.
    intro Heq.
    destruct f as [f_ob f_comm].
    destruct g as [g_ob g_comm].
    simpl in Heq.
    assert (Hob : f_ob = g_ob).
    {
      apply path_forall.
      exact Heq.
    }
    destruct Hob.
    f_ap.
    apply path_forall. intro n.
    apply path_ishprop.
  Qed.

  (* Composition of chain maps is associative *)
  Lemma comp_chain_map_assoc {A B C D : ChainComplex}
    (h : ChainMap C D) (g : ChainMap B C) (f : ChainMap A B) :
    comp_chain_map h (comp_chain_map g f) = comp_chain_map (comp_chain_map h g) f.
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply comp_hom_assoc.
  Qed.

  (* Composition with identity on the left *)
  Lemma comp_chain_map_id_left {A B : ChainComplex} (f : ChainMap A B) :
    comp_chain_map (id_chain_map B) f = f.
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply comp_hom_id_left.
  Qed.

  (* Composition with identity on the right *)
  Lemma comp_chain_map_id_right {A B : ChainComplex} (f : ChainMap A B) :
    comp_chain_map f (id_chain_map A) = f.
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply comp_hom_id_right.
  Qed.

  (* Helper: ChainMap forms a set *)
  Instance ChainMap_IsHSet `{Funext} (C D : ChainComplex) : IsHSet (ChainMap C D).
  Proof.
    (* ChainMap is equivalent to a sigma type *)
    assert (equiv_to_sig : ChainMap C D <~> 
      {f : forall n, GroupHom (ob C n) (ob D n) &
       forall n, comp_hom (f n) (diff C n) = comp_hom (diff D n) (f (S n))}).
    {
      apply (equiv_adjointify
        (fun cm => (map_ob C D cm; map_commutes C D cm))
        (fun p => Build_ChainMap C D p.1 p.2)).
      - (* Section *)
        intros [f Hf].
        reflexivity.
      - (* Retraction *)
        intros [f Hf].
        reflexivity.
    }
    (* Use the equivalence *)
    apply (istrunc_equiv_istrunc _ equiv_to_sig^-1).
  Qed.

  (* The category of chain complexes *)
  Definition ChainComplexCat `{Funext} : PreCategory.
  Proof.
    simple refine (@Build_PreCategory
      ChainComplex
      ChainMap
      id_chain_map
      (fun A B C => comp_chain_map)
      _ _ _ _).
    - (* associativity *)
      intros A B C D f g h.
      unfold comp_chain_map.
      apply ChainMap_eq.
      intro n.
      simpl.
      symmetry.
      apply comp_hom_assoc.
    - (* left identity *)
      intros A B f.
      apply comp_chain_map_id_left.
    - (* right identity *)
      intros A B f.
      apply comp_chain_map_id_right.
  Defined.

  (* The shift functor on chain complexes *)
  Definition ShiftComplex (C : ChainComplex) : ChainComplex.
  Proof.
    refine (Build_ChainComplex
      (fun n => ob C (S n))
      (fun n => diff C (S n))
      _).
    intro n.
    apply (diff_squared C (S n)).
  Defined.

  (* The shift functor on chain maps *)
  Definition ShiftMap {C D : ChainComplex} (f : ChainMap C D) : ChainMap (ShiftComplex C) (ShiftComplex D).
  Proof.
    refine (Build_ChainMap (ShiftComplex C) (ShiftComplex D)
      (fun n => map_ob C D f (S n))
      _).
    intro n.
    simpl.
    apply (map_commutes C D f (S n)).
  Defined.

  (* Helper: Composition with zero homomorphism is zero *)
  Lemma comp_zero_hom_left {A B C : AbelianGroupWithLaws} (f : GroupHom A B) :
    comp_hom (zero_hom B C) f = zero_hom A C.
  Proof.
    apply GroupHom_eq.
    reflexivity.
  Qed.

  (* Helper: Composition with zero homomorphism on the right is zero *)
  Lemma comp_zero_hom_right {A B C : AbelianGroupWithLaws} (f : GroupHom B C) :
    comp_hom f (zero_hom A B) = zero_hom A C.
  Proof.
    apply GroupHom_eq.
    apply path_forall. intro a.
    simpl.
    apply (hom_zero B C f).
  Qed.

  (* Replace the existing DesuspComplex definition *)
  Definition DesuspComplex (C : ChainComplex) : ChainComplex.
  Proof.
    simple refine (Build_ChainComplex _ _ _).
    - (* Objects: shift indices down by 1, with TrivialGroup at degree 0 *)
      intro n.
      destruct n as [|n'].
      + (* n = 0: We need something at degree 0 *)
        exact TrivialGroup.
      + (* n = S n': Use C at degree n' *)
        exact (ob C n').
    - (* Differential *)
      intro n.
      destruct n as [|n'].
      + (* d_0 : (DesuspComplex C)_1 → (DesuspComplex C)_0 
           That is: C_0 → TrivialGroup *)
        simpl.
        exact (zero_hom (ob C 0) TrivialGroup).
      + (* d_{n'+1} : C_{n'} → (previous degree) *)
        destruct n' as [|n''].
        * (* n' = 0, so we have d_1 : C_1 → C_0 *)
          simpl.
          exact (diff C 0).
        * (* n' = S n'', so we have d_{S(S n'')} : C_{S n''} → C_{n''} *)
          simpl.
          exact (diff C (S n'')).
    - (* Proof of diff_squared *)
      intro n.
      destruct n as [|n'].
      + (* n = 0: d_0 ∘ d_1 : C_1 → TrivialGroup *)
        simpl.
        (* d_0 is zero_hom, so composition with it is zero *)
        apply comp_zero_hom_left.
      + (* n = S n' *)
        destruct n' as [|n''].
        * (* n' = 0: d_1 ∘ d_2 *)
          simpl.
          apply (diff_squared C 0).
        * (* n' = S n'' *)
          simpl.
          apply (diff_squared C (S n'')).
  Defined.

  (* Replace the existing DesuspMap definition *)
  Definition DesuspMap {C D : ChainComplex} (f : ChainMap C D) : ChainMap (DesuspComplex C) (DesuspComplex D).
  Proof.
    simple refine (Build_ChainMap (DesuspComplex C) (DesuspComplex D) _ _).
    - (* map at each degree *)
      intro n.
      destruct n as [|n'].
      + (* n = 0: TrivialGroup → TrivialGroup *)
        simpl.
        exact (id_hom TrivialGroup).
      + (* n = S n': C_{n'} → D_{n'} *)
        simpl.
        exact (map_ob C D f n').
    - (* commutes with differential *)
      intro n.
      destruct n as [|n'].
      + (* n = 0: need to show 
           id ∘ zero_hom (ob C 0) TrivialGroup = zero_hom (ob D 0) TrivialGroup ∘ f_0 *)
        simpl.
        rewrite comp_hom_id_left.
        symmetry.
        apply comp_zero_hom_left.
      + (* n = S n' *)
        destruct n' as [|n''].
        * (* n' = 0 *)
          simpl.
          apply (map_commutes C D f 0).
        * (* n' = S n'' *)
          simpl.
          apply (map_commutes C D f (S n'')).
  Defined.

  (* Replace the existing epsilon_component definition *)
  Definition epsilon_component (C : ChainComplex) : ChainMap ((ShiftComplex o DesuspComplex) C) C.
  Proof.
    simpl.
    simple refine (Build_ChainMap (ShiftComplex (DesuspComplex C)) C _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      (* (Shift(Desusp(C)))_n = (Desusp(C))_{S n} = C_n *)
      exact (id_hom (ob C n)).
    - (* commutes with differential *)
      intro n.
      simpl.
      destruct n as [|n'].
      + (* n = 0 *)
        simpl.
        rewrite comp_hom_id_left.
        rewrite comp_hom_id_right.
        reflexivity.
      + (* n = S n' *)
        simpl.
        rewrite comp_hom_id_left.
        rewrite comp_hom_id_right.
        reflexivity.
  Defined.

  (* Replace the existing eta_component definition *)
  Definition eta_component (C : ChainComplex) : ChainMap C ((DesuspComplex o ShiftComplex) C).
  Proof.
    simpl.
    simple refine (Build_ChainMap C (DesuspComplex (ShiftComplex C)) _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      destruct n as [|n'].
      + (* n = 0: C_0 → TrivialGroup *)
        exact (zero_hom (ob C 0) TrivialGroup).
      + (* n = S n': C_{S n'} → (ShiftComplex C)_{n'} = C_{n'+1} = C_{S n'} *)
        exact (id_hom (ob C (S n'))).
    - (* commutes with differential *)
      intro n.
      destruct n as [|n'].
      + (* n = 0: need to show diff ∘ zero = zero ∘ diff *)
        simpl.
        rewrite comp_zero_hom_left.
        symmetry.
        rewrite comp_hom_id_right.
        reflexivity.
      + (* n = S n' *)
        destruct n' as [|n''].
        * (* n' = 0 *)
          simpl.
          rewrite comp_hom_id_left.
          rewrite comp_hom_id_right.
          reflexivity.
        * (* n' = S n'' *)
          simpl.
          rewrite comp_hom_id_left.
          rewrite comp_hom_id_right.
          reflexivity.
  Defined.

  (* Replace the existing eta_natural lemma *)
  Lemma eta_natural {C D : ChainComplex} (f : ChainMap C D) :
    comp_chain_map (DesuspMap (ShiftMap f)) (eta_component C) = 
    comp_chain_map (eta_component D) f.
  Proof.
    apply ChainMap_eq.
    intro n.
    destruct n as [|n'].
    - (* n = 0 *)
      simpl.
      apply GroupHom_eq.
      apply path_forall. intro a.
      simpl.
      (* Both sides are tt in TrivialGroup *)
      reflexivity.
    - (* n = S n' *)
      simpl.
      apply GroupHom_eq.
      apply path_forall. intro a.
      simpl.
      reflexivity.
  Qed.

  (* Replace the existing epsilon_natural lemma *)
  Lemma epsilon_natural {C D : ChainComplex} (f : ChainMap C D) :
    comp_chain_map f (epsilon_component C) = 
    comp_chain_map (epsilon_component D) (ShiftMap (DesuspMap f)).
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    destruct n as [|n'].
    - (* n = 0 *)
      simpl.
      reflexivity.
    - (* n = S n' *)
      simpl.
      reflexivity.
  Qed.

  (* Triangle identity 1: ε(Shift C) ∘ Shift(η C) = id on Shift C *)
  Lemma triangle_identity_1 (C : ChainComplex) :
    comp_chain_map (epsilon_component (ShiftComplex C)) (ShiftMap (eta_component C)) = 
    id_chain_map (ShiftComplex C).
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro a.
    simpl.
    reflexivity.
  Qed.

  (* Triangle identity 2: Desusp(ε C) ∘ η(Desusp C) = id on Desusp C *)
  Lemma triangle_identity_2 (C : ChainComplex) :
    comp_chain_map (DesuspMap (epsilon_component C)) (eta_component (DesuspComplex C)) = 
    id_chain_map (DesuspComplex C).
  Proof.
    apply ChainMap_eq.
    intro n.
    destruct n as [|n'].
    - (* n = 0 *)
      simpl.
      apply GroupHom_eq.
      apply path_forall. intro a.
      destruct a. (* a : Unit *)
      reflexivity.
    - (* n = S n' *)
      simpl.
      apply GroupHom_eq.
      apply path_forall. intro a.
      simpl.
      reflexivity.
  Qed.

  (* Make Desusp into a functor on ChainComplexCat *)
  Definition DesuspFunctor `{Funext} : Functor ChainComplexCat ChainComplexCat.
  Proof.
    refine (Build_Functor 
      ChainComplexCat ChainComplexCat
      DesuspComplex
      (fun C D => DesuspMap)
      _ _).
    - (* Functoriality: F(g ∘ f) = F(g) ∘ F(f) *)
      intros C D E f g.
      apply ChainMap_eq.
      intro n.
      destruct n as [|n'].
      + (* n = 0 *)
        simpl.
        reflexivity.
      + (* n = S n' *)
        simpl.
        reflexivity.
    - (* Preserves identity *)
      intro C.
      apply ChainMap_eq.
      intro n.
      destruct n as [|n'].
      + (* n = 0 *)
        simpl.
        reflexivity.
      + (* n = S n' *)
        simpl.
        reflexivity.
  Defined.

  (* Make Shift into a functor on ChainComplexCat *)
  Definition ShiftFunctor `{Funext} : Functor ChainComplexCat ChainComplexCat.
  Proof.
    refine (Build_Functor 
      ChainComplexCat ChainComplexCat
      ShiftComplex
      (fun C D => ShiftMap)
      _ _).
    - (* Functoriality: F(g ∘ f) = F(g) ∘ F(f) *)
      intros C D E f g.
      apply ChainMap_eq.
      intro n.
      reflexivity.
    - (* Preserves identity *)
      intro C.
      apply ChainMap_eq.
      intro n.
      reflexivity.
  Defined.

  (* Create the unit natural transformation η : Id → Desusp ∘ Shift *)
  Definition eta_chain `{Funext} : NaturalTransformation 
    (1%functor : Functor ChainComplexCat ChainComplexCat)
    ((DesuspFunctor o ShiftFunctor)%functor).
  Proof.
    refine (Build_NaturalTransformation _ _ 
      (fun C => eta_component C : morphism ChainComplexCat 
                                    (object_of 1%functor C)
                                    (object_of (DesuspFunctor o ShiftFunctor)%functor C)) _).
    intros C D f.
    simpl.
    symmetry.
    exact (eta_natural f).
  Defined.

  (* Create the counit natural transformation ε : Shift ∘ Desusp → Id *)
  Definition epsilon_chain `{Funext} : NaturalTransformation 
    ((ShiftFunctor o DesuspFunctor)%functor)
    (1%functor : Functor ChainComplexCat ChainComplexCat).
  Proof.
    refine (Build_NaturalTransformation _ _ 
      (fun C => epsilon_component C : morphism ChainComplexCat 
                                        (object_of (ShiftFunctor o DesuspFunctor)%functor C)
                                        (object_of 1%functor C)) _).
    intros C D f.
    simpl.
    symmetry.
    exact (epsilon_natural f).
  Defined.

  Definition ZeroChainComplex : ChainComplex.
  Proof.
    refine (Build_ChainComplex
      (fun n => TrivialGroup)
      (fun n => zero_hom TrivialGroup TrivialGroup)
      _).
    intro n.
    apply comp_zero_hom_left.
  Defined.

  Definition DirectSumChainComplex (C D : ChainComplex) : ChainComplex.
  Proof.
    simple refine (Build_ChainComplex
      (fun n => DirectSum (ob C n) (ob D n))
      _ _).
    - (* differential *)
      intro n.
      simple refine (Build_GroupHom _ _ _ _ _).
      + (* map *)
        exact (fun p => (hom_map _ _ (diff C n) (fst p), 
                         hom_map _ _ (diff D n) (snd p))).
      + (* hom_zero *)
        simpl.
        f_ap.
        * apply (hom_zero _ _ (diff C n)).
        * apply (hom_zero _ _ (diff D n)).
      + (* hom_plus *)
        intros [c1 d1] [c2 d2].
        simpl.
        f_ap.
        * apply (hom_plus _ _ (diff C n)).
        * apply (hom_plus _ _ (diff D n)).
    - (* diff_squared *)
      intro n.
      apply GroupHom_eq.
      apply path_forall. intro p.
      destruct p as [c d].
      simpl.
      pose proof (diff_squared C n) as HC.
      pose proof (diff_squared D n) as HD.
      pose proof (ap (fun h => hom_map _ _ h c) HC) as Hc.
      pose proof (ap (fun h => hom_map _ _ h d) HD) as Hd.
      simpl in Hc, Hd.
      f_ap; assumption.
  Defined.

  Theorem ZeroChainComplex_is_zero : ZeroObject ChainComplexCat.
  Proof.
    refine (Build_ZeroObject ChainComplexCat ZeroChainComplex _ _).
    - (* initial *)
      intro C.
      simple refine (Build_Contr _ _ _).
      + (* center: the zero chain map *)
        simple refine (Build_ChainMap ZeroChainComplex C _ _).
        * (* map at each degree *)
          intro n.
          apply zero_hom.
        * (* commutes *)
          intro n.
          simpl.
          rewrite comp_zero_hom_left.
          rewrite comp_zero_hom_right.
          reflexivity.
      + (* contr *)
        intro f.
        apply ChainMap_eq.
        intro n.
        apply GroupHom_eq.
        apply path_forall. intro x.
        destruct x.
        simpl.
        symmetry.
        exact (hom_zero _ _ (map_ob _ _ f n)).
    - (* terminal *)
      intro C.
      simple refine (Build_Contr _ _ _).
      + (* center *)
        simple refine (Build_ChainMap C ZeroChainComplex _ _).
        * (* map at each degree *)
          intro n.
          apply zero_hom.
        * (* commutes *)
          intro n.
          simpl.
          rewrite comp_zero_hom_left.
          rewrite comp_zero_hom_right.
          reflexivity.
      + (* contr *)
        intro f.
        apply ChainMap_eq.
        intro n.
        apply GroupHom_eq.
        apply path_forall. intro x.
        destruct (hom_map _ _ (map_ob _ _ f n) x).
        reflexivity.
  Defined.

  Definition chain_inj1 (C D : ChainComplex) : ChainMap C (DirectSumChainComplex C D).
  Proof.
    simple refine (Build_ChainMap C (DirectSumChainComplex C D) _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      exact (inj1 (ob C n) (ob D n)).
    - (* commutes *)
      intro n.
      apply GroupHom_eq.
      apply path_forall. intro c.
      simpl.
      f_ap.
      symmetry.
      apply (hom_zero _ _ (diff D n)).
  Defined.

  Definition chain_inj2 (C D : ChainComplex) : ChainMap D (DirectSumChainComplex C D).
  Proof.
    simple refine (Build_ChainMap D (DirectSumChainComplex C D) _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      exact (inj2 (ob C n) (ob D n)).
    - (* commutes *)
      intro n.
      apply GroupHom_eq.
      apply path_forall. intro d.
      simpl.
      f_ap.
      symmetry.
      apply (hom_zero _ _ (diff C n)).
  Defined.

  Definition chain_proj1 (C D : ChainComplex) : ChainMap (DirectSumChainComplex C D) C.
  Proof.
    simple refine (Build_ChainMap (DirectSumChainComplex C D) C _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      exact (proj1 (ob C n) (ob D n)).
    - (* commutes *)
      intro n.
      apply GroupHom_eq.
      apply path_forall. intros [c d].
      reflexivity.
  Defined.

  Definition chain_proj2 (C D : ChainComplex) : ChainMap (DirectSumChainComplex C D) D.
  Proof.
    simple refine (Build_ChainMap (DirectSumChainComplex C D) D _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      exact (proj2 (ob C n) (ob D n)).
    - (* commutes *)
      intro n.
      apply GroupHom_eq.
      apply path_forall. intros [c d].
      reflexivity.
  Defined.

  Lemma chain_beta_l (C D : ChainComplex) : 
    comp_chain_map (chain_proj1 C D) (chain_inj1 C D) = id_chain_map C.
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro c.
    reflexivity.
  Qed.

  Lemma chain_beta_r (C D : ChainComplex) : 
    comp_chain_map (chain_proj2 C D) (chain_inj2 C D) = id_chain_map D.
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro d.
    reflexivity.
  Qed.

  Definition zero_chain_map (C D : ChainComplex) : ChainMap C D.
  Proof.
    simple refine (Build_ChainMap C D _ _).
    - (* map at each degree *)
      intro n.
      apply zero_hom.
    - (* commutes *)
      intro n.
      rewrite comp_zero_hom_left.
      rewrite comp_zero_hom_right.
      reflexivity.
  Defined.

  Lemma chain_mixed_l (C D : ChainComplex) : 
    comp_chain_map (chain_proj1 C D) (chain_inj2 C D) = zero_chain_map D C.
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro d.
    reflexivity.
  Qed.

  Lemma chain_mixed_r (C D : ChainComplex) : 
    comp_chain_map (chain_proj2 C D) (chain_inj1 C D) = zero_chain_map C D.
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro c.
    reflexivity.
  Qed.

  Lemma zero_chain_map_is_zero_morphism (C D : ChainComplex) :
    zero_chain_map C D = zero_morphism ZeroChainComplex_is_zero C D.
  Proof.
    unfold zero_morphism.
    simpl.
    apply ChainMap_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intro c.
    simpl.
    reflexivity.
  Qed.

  Definition chain_coprod_mor (C D W : ChainComplex) 
    (f : ChainMap C W) (g : ChainMap D W) : ChainMap (DirectSumChainComplex C D) W.
  Proof.
    simple refine (Build_ChainMap (DirectSumChainComplex C D) W _ _).
    - (* map at each degree *)
      intro n.
      simple refine (Build_GroupHom _ _ _ _ _).
      + (* map *)
        intros [c d].
        exact (plus (group (ob W n))
          (hom_map _ _ (map_ob C W f n) c)
          (hom_map _ _ (map_ob D W g n) d)).
      + (* hom_zero *)
        simpl.
        rewrite (hom_zero _ _ (map_ob C W f n)).
        rewrite (hom_zero _ _ (map_ob D W g n)).
        apply (plus_zero_l _ (laws (ob W n))).
      + (* hom_plus *)
        intros [c1 d1] [c2 d2].
        simpl.
        rewrite (hom_plus _ _ (map_ob C W f n)).
        rewrite (hom_plus _ _ (map_ob D W g n)).
        (* Goal: (f c1 + g d1) + (f c2 + g d2) = (f c1 + f c2) + (g d1 + g d2) *)
        set (fc1 := hom_map _ _ (map_ob C W f n) c1).
        set (fc2 := hom_map _ _ (map_ob C W f n) c2).
        set (gd1 := hom_map _ _ (map_ob D W g n) d1).
        set (gd2 := hom_map _ _ (map_ob D W g n) d2).
        (* Apply associativity and commutativity *)
        rewrite <- (plus_assoc _ (laws (ob W n)) fc1 gd1 _).
        rewrite (plus_assoc _ (laws (ob W n)) gd1 fc2 gd2).
        rewrite (plus_comm _ (laws (ob W n)) gd1 fc2).
        rewrite <- (plus_assoc _ (laws (ob W n)) fc2 gd1 gd2).
        rewrite (plus_assoc _ (laws (ob W n)) fc1 fc2 _).
        reflexivity.
    - (* commutes *)
      intro n.
      apply GroupHom_eq.
      apply path_forall. intros [c d].
      simpl.
      pose proof (map_commutes C W f n) as Hf.
      pose proof (map_commutes D W g n) as Hg.
      apply (ap (fun h => hom_map _ _ h c)) in Hf.
      apply (ap (fun h => hom_map _ _ h d)) in Hg.
      simpl in Hf, Hg.
      rewrite Hf, Hg.
      symmetry.
      apply (hom_plus _ _ (diff W n)).
  Defined.

  Lemma chain_coprod_beta_l (C D W : ChainComplex) 
    (f : ChainMap C W) (g : ChainMap D W) :
    comp_chain_map (chain_coprod_mor C D W f g) (chain_inj1 C D) = f.
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro c.
    simpl.
    rewrite (hom_zero _ _ (map_ob D W g n)).
    apply (plus_zero_r _ (laws (ob W n))).
  Qed.

  Lemma chain_coprod_beta_r (C D W : ChainComplex) 
    (f : ChainMap C W) (g : ChainMap D W) :
    comp_chain_map (chain_coprod_mor C D W f g) (chain_inj2 C D) = g.
  Proof.
    apply ChainMap_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro d.
    simpl.
    rewrite (hom_zero _ _ (map_ob C W f n)).
    apply (plus_zero_l _ (laws (ob W n))).
  Qed.

  Lemma chain_coprod_unique (C D W : ChainComplex) 
    (f : ChainMap C W) (g : ChainMap D W)
    (h : ChainMap (DirectSumChainComplex C D) W) :
    comp_chain_map h (chain_inj1 C D) = f ->
    comp_chain_map h (chain_inj2 C D) = g ->
    h = chain_coprod_mor C D W f g.
  Proof.
    intros Hf Hg.
    apply ChainMap_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intros [c d].
    (* Express (c,d) as a sum in DirectSum *)
    assert (Heq : (c, d) = plus (group (DirectSum (ob C n) (ob D n)))
                                 (c, zero (group (ob D n))) 
                                 (zero (group (ob C n)), d)).
    {
      simpl.
      f_ap.
      - symmetry. apply (plus_zero_r _ (laws (ob C n))).
      - symmetry. apply (plus_zero_l _ (laws (ob D n))).
    }
    rewrite Heq.
    rewrite (hom_plus _ _ (map_ob _ _ h n)).
    (* Use the fact that h ∘ inj1 = f at degree n *)
    assert (Hfc : hom_map _ _ (map_ob _ _ h n) (c, zero (group (ob D n))) = 
                  hom_map _ _ (map_ob C W f n) c).
    {
      change (hom_map _ _ (map_ob _ _ h n) (hom_map _ _ (inj1 _ _) c) = 
              hom_map _ _ (map_ob C W f n) c).
      unfold comp_hom.
      pose proof (ap (fun k => map_ob _ _ k n) Hf) as Hf_n.
      exact (ap (fun k => hom_map _ _ k c) Hf_n).
    }
    (* Use the fact that h ∘ inj2 = g at degree n *)
    assert (Hgd : hom_map _ _ (map_ob _ _ h n) (zero (group (ob C n)), d) = 
                  hom_map _ _ (map_ob D W g n) d).
    {
      change (hom_map _ _ (map_ob _ _ h n) (hom_map _ _ (inj2 _ _) d) = 
              hom_map _ _ (map_ob D W g n) d).
      unfold comp_hom.
      pose proof (ap (fun k => map_ob _ _ k n) Hg) as Hg_n.
      exact (ap (fun k => hom_map _ _ k d) Hg_n).
    }
    rewrite Hfc, Hgd.
    (* Now simplify the goal *)
    simpl.
    (* Need to handle the extra plus terms *)
    rewrite (plus_zero_r _ (laws (ob C n))).
    rewrite (plus_zero_l _ (laws (ob D n))).
    reflexivity.
  Qed.

  Definition chain_prod_mor (W C D : ChainComplex) 
    (f : ChainMap W C) (g : ChainMap W D) : ChainMap W (DirectSumChainComplex C D).
  Proof.
    simple refine (Build_ChainMap W (DirectSumChainComplex C D) _ _).
    - (* map at each degree *)
      intro n.
      simple refine (Build_GroupHom _ _ _ _ _).
      + (* map *)
        intro w.
        exact (hom_map _ _ (map_ob W C f n) w,
               hom_map _ _ (map_ob W D g n) w).
      + (* hom_zero *)
        simpl.
        f_ap.
        * apply (hom_zero _ _ (map_ob W C f n)).
        * apply (hom_zero _ _ (map_ob W D g n)).
      + (* hom_plus *)
        intros w1 w2.
        simpl.
        f_ap.
        * apply (hom_plus _ _ (map_ob W C f n)).
        * apply (hom_plus _ _ (map_ob W D g n)).
    - (* commutes *)
      intro n.
      apply GroupHom_eq.
      apply path_forall. intro w.
      simpl.
      pose proof (map_commutes W C f n) as Hf.
      pose proof (map_commutes W D g n) as Hg.
      apply (ap (fun h => hom_map _ _ h w)) in Hf.
      apply (ap (fun h => hom_map _ _ h w)) in Hg.
      simpl in Hf, Hg.
      f_ap; assumption.
  Defined.

  Lemma chain_prod_beta_l (W C D : ChainComplex) 
    (f : ChainMap W C) (g : ChainMap W D) :
    comp_chain_map (chain_proj1 C D) (chain_prod_mor W C D f g) = f.
  Proof.
    apply ChainMap_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intro w.
    reflexivity.
  Qed.

  Lemma chain_prod_beta_r (W C D : ChainComplex) 
    (f : ChainMap W C) (g : ChainMap W D) :
    comp_chain_map (chain_proj2 C D) (chain_prod_mor W C D f g) = g.
  Proof.
    apply ChainMap_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intro w.
    reflexivity.
  Qed.

  Lemma chain_prod_unique (W C D : ChainComplex) 
    (f : ChainMap W C) (g : ChainMap W D)
    (h : ChainMap W (DirectSumChainComplex C D)) :
    comp_chain_map (chain_proj1 C D) h = f ->
    comp_chain_map (chain_proj2 C D) h = g ->
    h = chain_prod_mor W C D f g.
  Proof.
    intros Hf Hg.
    apply ChainMap_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intro w.
    pose proof (ap (fun k => map_ob _ _ k n) Hf) as Hf_n.
    pose proof (ap (fun k => map_ob _ _ k n) Hg) as Hg_n.
    pose proof (ap (fun k => hom_map _ _ k w) Hf_n) as Hc.
    pose proof (ap (fun k => hom_map _ _ k w) Hg_n) as Hd.
    simpl in Hc, Hd.
    destruct (hom_map _ _ (map_ob _ _ h n) w) as [c d].
    simpl in *.
    f_ap; assumption.
  Qed.

  Definition ChainComplexBiproduct (C D : ChainComplex) : @Biproduct ChainComplexCat C D ZeroChainComplex_is_zero.
  Proof.
    (* Biproduct data *)
    pose (bdata := Build_BiproductData ChainComplexCat C D 
      (DirectSumChainComplex C D)
      (chain_inj1 C D)
      (chain_inj2 C D)
      (chain_proj1 C D)
      (chain_proj2 C D)).
      
    (* Biproduct axioms *)
    assert (bis : IsBiproduct bdata ZeroChainComplex_is_zero).
    {
      simple refine (Build_IsBiproduct _ _ _ _ _ _ _ _ _).
      - apply chain_beta_l.
      - apply chain_beta_r.
      - rewrite <- zero_chain_map_is_zero_morphism. apply chain_mixed_l.
      - rewrite <- zero_chain_map_is_zero_morphism. apply chain_mixed_r.
    }
    
    (* Universal property *)
    assert (buni : HasBiproductUniversal bdata).
    {
      simple refine (Build_HasBiproductUniversal _ _ _ _ _ _).
      - (* Coproduct universal *)
        intros W f g.
        apply (Build_Contr _ (chain_coprod_mor C D W f g; (chain_coprod_beta_l C D W f g, chain_coprod_beta_r C D W f g))).
        intros [h [Hl Hr]].
        simpl.
        apply path_sigma_uncurried.
        simpl.
        exists ((chain_coprod_unique C D W f g h Hl Hr)^).
        apply path_ishprop.
      - (* Product universal *)
        intros W f g.
        apply (Build_Contr _ (chain_prod_mor W C D f g; (chain_prod_beta_l W C D f g, chain_prod_beta_r W C D f g))).
        intros [h [Hl Hr]].
        simpl.
        apply path_sigma_uncurried.
        simpl.
        exists ((chain_prod_unique W C D f g h Hl Hr)^).
        apply path_ishprop.
    }
    
    exact (Build_Biproduct _ _ _ _ bdata bis buni).
  Defined.

  Definition ChainComplexAdditive `{Funext} : AdditiveCategory.
  Proof.
    exact (Build_AdditiveCategory 
      ChainComplexCat
      ZeroChainComplex_is_zero
      ChainComplexBiproduct).
  Defined.

  Definition shift_zero_iso : ChainMap (ShiftComplex ZeroChainComplex) ZeroChainComplex.
  Proof.
    simple refine (Build_ChainMap _ _ _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      exact (id_hom TrivialGroup).
    - (* commutes *)
      intro n.
      simpl.
      reflexivity.
  Defined.

  Definition shift_zero_iso_inv : ChainMap ZeroChainComplex (ShiftComplex ZeroChainComplex).
  Proof.
    simple refine (Build_ChainMap _ _ _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      exact (id_hom TrivialGroup).
    - (* commutes *)
      intro n.
      simpl.
      reflexivity.
  Defined.

  Lemma ShiftFunctor_preserves_zero_iso : 
    comp_chain_map shift_zero_iso shift_zero_iso_inv = id_chain_map ZeroChainComplex /\
    comp_chain_map shift_zero_iso_inv shift_zero_iso = id_chain_map (ShiftComplex ZeroChainComplex).
  Proof.
    split.
    - apply ChainMap_eq. intro n. simpl. reflexivity.
    - apply ChainMap_eq. intro n. simpl. reflexivity.
  Qed.

  Definition shift_biproduct_iso (C D : ChainComplex) : 
    ChainMap (ShiftComplex (DirectSumChainComplex C D)) 
             (DirectSumChainComplex (ShiftComplex C) (ShiftComplex D)).
  Proof.
    simple refine (Build_ChainMap _ _ _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      exact (id_hom (DirectSum (ob C (S n)) (ob D (S n)))).
    - (* commutes *)
      intro n.
      simpl.
      reflexivity.
  Defined.

  Definition shift_biproduct_iso_inv (C D : ChainComplex) : 
    ChainMap (DirectSumChainComplex (ShiftComplex C) (ShiftComplex D))
             (ShiftComplex (DirectSumChainComplex C D)).
  Proof.
    simple refine (Build_ChainMap _ _ _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      exact (id_hom (DirectSum (ob C (S n)) (ob D (S n)))).
    - (* commutes *)
      intro n.
      simpl.
      reflexivity.
  Defined.

  Lemma shift_biproduct_iso_is_iso (C D : ChainComplex) :
    comp_chain_map (shift_biproduct_iso C D) (shift_biproduct_iso_inv C D) = 
    id_chain_map (DirectSumChainComplex (ShiftComplex C) (ShiftComplex D)) /\
    comp_chain_map (shift_biproduct_iso_inv C D) (shift_biproduct_iso C D) = 
    id_chain_map (ShiftComplex (DirectSumChainComplex C D)).
  Proof.
    split.
    - apply ChainMap_eq. intro n. simpl. reflexivity.
    - apply ChainMap_eq. intro n. simpl. reflexivity.
  Qed.


  (* Desusp preserves the zero object *)
  Definition desusp_zero_iso : ChainMap (DesuspComplex ZeroChainComplex) ZeroChainComplex.
  Proof.
    simple refine (Build_ChainMap _ _ _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      destruct n as [|n'].
      + (* n = 0: TrivialGroup → TrivialGroup *)
        exact (id_hom TrivialGroup).
      + (* n = S n': TrivialGroup → TrivialGroup *)
        exact (id_hom TrivialGroup).
    - (* commutes *)
      intro n.
      simpl.
      destruct n as [|n'].
      + (* n = 0 *)
        simpl.
        reflexivity.
      + (* n = S n' *)
        destruct n' as [|n''].
        * (* n' = 0 *)
          simpl.
          reflexivity.
        * (* n' = S n'' *)
          simpl.
          reflexivity.
  Defined.

  Definition desusp_zero_iso_inv : ChainMap ZeroChainComplex (DesuspComplex ZeroChainComplex).
  Proof.
    simple refine (Build_ChainMap _ _ _ _).
    - (* map at each degree *)
      intro n.
      simpl.
      destruct n as [|n'].
      + (* n = 0: TrivialGroup → TrivialGroup *)
        exact (id_hom TrivialGroup).
      + (* n = S n': TrivialGroup → TrivialGroup *)
        exact (id_hom TrivialGroup).
    - (* commutes *)
      intro n.
      simpl.
      destruct n as [|n'].
      + (* n = 0 *)
        simpl.
        reflexivity.
      + (* n = S n' *)
        destruct n' as [|n''].
        * (* n' = 0 *)
          simpl.
          reflexivity.
        * (* n' = S n'' *)
          simpl.
          reflexivity.
  Defined.

  Lemma DesuspFunctor_preserves_zero_iso : 
    comp_chain_map desusp_zero_iso desusp_zero_iso_inv = id_chain_map ZeroChainComplex /\
    comp_chain_map desusp_zero_iso_inv desusp_zero_iso = id_chain_map (DesuspComplex ZeroChainComplex).
  Proof.
    split.
    - (* First part: desusp_zero_iso ∘ desusp_zero_iso_inv = id on ZeroChainComplex *)
      apply ChainMap_eq. 
      intro n.
      destruct n; reflexivity.
      
    - (* Second part: desusp_zero_iso_inv ∘ desusp_zero_iso = id on DesuspComplex ZeroChainComplex *)
      apply ChainMap_eq. 
      intro n.
      destruct n; reflexivity.
  Qed.

  (* Shift is an additive functor *)
  Definition ShiftAdditiveFunctor `{Funext} : AdditiveFunctor ChainComplexAdditive ChainComplexAdditive.
  Proof.
    refine (Build_AdditiveFunctor 
      ChainComplexAdditive ChainComplexAdditive
      ShiftFunctor
      _ _).
    - (* preserves_zero *)
      simpl.
      (* ShiftComplex ZeroChainComplex = ZeroChainComplex up to isomorphism *)
      reflexivity.
    - (* preserves_biproduct *)
      intros C D.
      simpl.
      (* ShiftComplex (DirectSumChainComplex C D) = 
         DirectSumChainComplex (ShiftComplex C) (ShiftComplex D) *)
      reflexivity.
  Defined.

  Lemma desusp_zero_objects_eq (n : nat) : 
    ob (DesuspComplex ZeroChainComplex) n = ob ZeroChainComplex n.
  Proof.
    destruct n; reflexivity.
  Qed.

  (* Helper lemma: the object function simplifies correctly *)
  Lemma desusp_zero_ob_eq : 
    (fun n : nat => match n with | 0%nat => TrivialGroup | S _ => TrivialGroup end) = 
    (fun n : nat => TrivialGroup).
  Proof.
    apply path_forall. intro n.
    destruct n; reflexivity.
  Qed.

  (* Helper lemma: the differential function simplifies correctly *)
  Lemma desusp_zero_diff_eq :
    (fun n : nat => match n with 
                    | 0%nat => zero_hom TrivialGroup TrivialGroup
                    | S _ => zero_hom TrivialGroup TrivialGroup 
                    end) =
    (fun n : nat => zero_hom TrivialGroup TrivialGroup).
  Proof.
    apply path_forall. intro n.
    destruct n; reflexivity.
  Qed.

  Lemma ChainComplex_eq (C D : ChainComplex) 
    (Hob : ob C = ob D)
    (Hdiff : forall n, transport (fun ob_fun => GroupHom (ob_fun (S n)) (ob_fun n)) 
                                 Hob 
                                 (diff C n) = diff D n) :
    C = D.
  Proof.
    destruct C as [obC diffC sqC].
    destruct D as [obD diffD sqD].
    simpl in *.
    destruct Hob.
    simpl in Hdiff.
    assert (Hd : diffC = diffD).
    { apply path_forall. exact Hdiff. }
    destruct Hd.
    f_ap.
    apply path_forall. intro n.
    apply path_ishprop.
  Qed.

  Lemma desusp_zero_preserves : 
    DesuspComplex ZeroChainComplex = ZeroChainComplex.
  Proof.
    assert (ob_eq : ob (DesuspComplex ZeroChainComplex) = ob ZeroChainComplex).
    { apply path_forall. intro n. destruct n; reflexivity. }
    
    assert (diff_eq : forall n, 
      transport (fun f => GroupHom (f (S n)) (f n)) ob_eq 
                (diff (DesuspComplex ZeroChainComplex) n) = 
      diff ZeroChainComplex n).
    {
      intro n.
      (* Key insight: there's only one homomorphism TrivialGroup → TrivialGroup *)
      assert (unique_hom : forall (f g : GroupHom TrivialGroup TrivialGroup), f = g).
      {
        intros f g.
        apply GroupHom_eq.
        apply path_forall. intro x.
        destruct x. 
        destruct (hom_map _ _ f tt), (hom_map _ _ g tt).
        reflexivity.
      }
      (* Apply this to our transported morphism *)
      apply unique_hom.
    }
    
    exact (ChainComplex_eq _ _ ob_eq diff_eq).
  Qed.

  Definition trivial_to_directsum_trivial : 
    GroupHom TrivialGroup (DirectSum TrivialGroup TrivialGroup).
  Proof.
    refine (Build_GroupHom TrivialGroup (DirectSum TrivialGroup TrivialGroup) 
      (fun _ => (zero (group TrivialGroup), zero (group TrivialGroup))) _ _).
    - (* hom_zero *)
      reflexivity.
    - (* hom_plus *)
      intros x y. 
      simpl.
      destruct x, y.
      reflexivity.
  Defined.

  Definition desusp_biproduct_iso (C D : ChainComplex) : 
    ChainMap (DesuspComplex (DirectSumChainComplex C D))
             (DirectSumChainComplex (DesuspComplex C) (DesuspComplex D)).
  Proof.
    simple refine (Build_ChainMap _ _ _ _).
    - (* map at each degree *)
      intro n.
      destruct n as [|n'].
      + (* n = 0: TrivialGroup → DirectSum TrivialGroup TrivialGroup *)
        exact trivial_to_directsum_trivial.
      + (* n = S n': DirectSum (ob C n') (ob D n') → DirectSum (ob C n') (ob D n') *)
        exact (id_hom _).
    - (* commutes *)
      intro n.
      destruct n as [|n'].
      + (* n = 0 *)
        apply GroupHom_eq.
        apply path_forall. intro x.
        destruct x. reflexivity.
      + (* n = S n' *)
        destruct n' as [|n''].
        * (* n' = 0: special case where codomain changes *)
          simpl.
          apply GroupHom_eq.
          apply path_forall. intros [c d].
          simpl.
          reflexivity.
        * (* n' = S n'' *)
          simpl.
          (* Both differentials are the same, and composing with identity gives identity *)
          reflexivity.
  Defined.

  Definition desusp_biproduct_iso_inv (C D : ChainComplex) : 
    ChainMap (DirectSumChainComplex (DesuspComplex C) (DesuspComplex D))
             (DesuspComplex (DirectSumChainComplex C D)).
  Proof.
    simple refine (Build_ChainMap _ _ _ _).
    - (* map at each degree *)
      intro n.
      destruct n as [|n'].
      + (* n = 0: DirectSum TrivialGroup TrivialGroup → TrivialGroup *)
        exact (zero_hom _ _).
      + (* n = S n': DirectSum (ob C n') (ob D n') → DirectSum (ob C n') (ob D n') *)
        exact (id_hom _).
    - (* commutes *)
      intro n.
      destruct n as [|n'].
      + (* n = 0 *)
        simpl.
        rewrite comp_zero_hom_right.
        rewrite comp_zero_hom_left.
        reflexivity.
      + (* n = S n' *)
        destruct n' as [|n''].
        * (* n' = 0 *)
          simpl.
          reflexivity.
        * (* n' = S n'' *)
          simpl.
          reflexivity.
  Defined.

  Lemma desusp_biproduct_iso_is_iso (C D : ChainComplex) :
    comp_chain_map (desusp_biproduct_iso C D) (desusp_biproduct_iso_inv C D) = 
    id_chain_map (DirectSumChainComplex (DesuspComplex C) (DesuspComplex D)) /\
    comp_chain_map (desusp_biproduct_iso_inv C D) (desusp_biproduct_iso C D) = 
    id_chain_map (DesuspComplex (DirectSumChainComplex C D)).
  Proof.
    split.
    - (* First direction *)
      apply ChainMap_eq.
      intro n.
      destruct n as [|n'].
      + (* n = 0 *)
        simpl.
        apply GroupHom_eq.
        apply path_forall. intros [t1 t2].
        destruct t1, t2.
        reflexivity.
      + (* n = S n' *)
        simpl.
        reflexivity.
    - (* Second direction *)
      apply ChainMap_eq.
      intro n.
      destruct n as [|n'].
      + (* n = 0 *)
        simpl.
        apply GroupHom_eq.
        apply path_forall. intro t.
        destruct t.
        reflexivity.
      + (* n = S n' *)
        simpl.
        reflexivity.
  Qed.

  (* Define Loop functor differently to ensure it preserves biproducts *)
  Definition LoopComplex (C : ChainComplex) : ChainComplex.
  Proof.
    simple refine (Build_ChainComplex _ _ _).
    - (* Objects: insert TrivialGroup at degree 0, shift everything else up *)
      intro n.
      exact (ob C (S n)).
    - (* Differential *)
      intro n.
      exact (diff C (S n)).
    - (* diff_squared *)
      intro n.
      exact (diff_squared C (S n)).
  Defined.

  (** * A trivial pre-stable structure on TwoAdditive *)

  Definition TrivialSuspLoop : AdditiveFunctor TwoCatAdditive.TwoAdditive TwoCatAdditive.TwoAdditive.
  Proof.
    refine (Build_AdditiveFunctor 
      TwoCatAdditive.TwoAdditive TwoCatAdditive.TwoAdditive
      1%functor  (* identity functor *)
      _ _).
    - (* preserves_zero *)
      reflexivity.
    - (* preserves_biproduct *)
      intros X Y.
      reflexivity.
  Defined.

  Definition TrivialEta : NaturalTransformation 1%functor (TrivialSuspLoop o TrivialSuspLoop)%functor.
  Proof.
    refine (Build_NaturalTransformation _ _ 
      (fun X => 1%morphism) _).
    intros X Y f.
    simpl.
    (* id ∘ f = f ∘ id in TwoCat *)
    destruct X, Y; destruct f; reflexivity.
  Defined.

  Definition TrivialEpsilon : NaturalTransformation (TrivialSuspLoop o TrivialSuspLoop)%functor 1%functor.
  Proof.
    refine (Build_NaturalTransformation _ _ 
      (fun X => 1%morphism) _).
    intros X Y f.
    simpl.
    destruct X, Y; destruct f; reflexivity.
  Defined.

  Definition TrivialPreStable : PreStableCategory.
  Proof.
    exact (Build_PreStableCategory
      TwoCatAdditive.TwoAdditive
      TrivialSuspLoop
      TrivialSuspLoop
      TrivialEta
      TrivialEpsilon).
  Defined.

  Lemma two_id_left_identity (X Y : SimpleBiproductCategory.TwoObj) 
    (f : SimpleBiproductCategory.TwoMor X Y) :
    SimpleBiproductCategory.two_comp (SimpleBiproductCategory.two_id Y) f = f.
  Proof.
    destruct X, Y; destruct f; reflexivity.
  Qed.

  Lemma two_id_right_identity (X Y : SimpleBiproductCategory.TwoObj) 
    (f : SimpleBiproductCategory.TwoMor X Y) :
    SimpleBiproductCategory.two_comp f (SimpleBiproductCategory.two_id X) = f.
  Proof.
    destruct X, Y; destruct f; reflexivity.
  Qed.

  Lemma two_id_is_identity (X : SimpleBiproductCategory.TwoObj) :
    @SimpleBiproductCategory.two_id X = @Category.Core.identity SimpleBiproductCategory.TwoCat X.
  Proof.
    destruct X; reflexivity.
  Qed.

  Definition id_morphism_is_iso (C : PreCategory) (X : C) :
    IsIsomorphism (1%morphism : morphism C X X).
  Proof.
    exact (Build_IsIsomorphism C X X 1%morphism 1%morphism 
             (left_identity C X X 1%morphism)
             (right_identity C X X 1%morphism)).
  Defined.

  Lemma TrivialEta_is_iso : forall X, IsIsomorphism (components_of TrivialEta X).
  Proof.
    intro X.
    simpl.
    apply id_morphism_is_iso.
  Qed.

  Lemma TrivialEpsilon_is_iso : forall X, IsIsomorphism (components_of TrivialEpsilon X).
  Proof.
    intro X.
    simpl.
    apply id_morphism_is_iso.
  Qed.

  Lemma TrivialTriangle1 : forall X,
    (components_of TrivialEpsilon (object_of TrivialSuspLoop X) o 
     morphism_of TrivialSuspLoop (components_of TrivialEta X))%morphism = 1%morphism.
  Proof.
    intro X.
    simpl.
    apply two_id_left_identity.
  Qed.

  Lemma TrivialTriangle2 : forall X,
    (morphism_of TrivialSuspLoop (components_of TrivialEpsilon X) o
     components_of TrivialEta (object_of TrivialSuspLoop X))%morphism = 1%morphism.
  Proof.
    intro X.
    simpl.
    apply two_id_left_identity.
  Qed.

  Require Import ProperStableCategories.

  Lemma TrivialEta_is_iso_proper : forall X, 
    OppositeCategories.IsIsomorphism (components_of (eta TrivialPreStable) X).
  Proof.
    intro X.
    simpl.
    exists 1%morphism.
    split.
    - apply two_id_left_identity.
    - apply two_id_right_identity.
  Qed.

  Lemma TrivialEpsilon_is_iso_proper : forall X, 
    OppositeCategories.IsIsomorphism (components_of (epsilon TrivialPreStable) X).
  Proof.
    intro X.
    simpl.
    exists 1%morphism.
    split.
    - apply two_id_left_identity.
    - apply two_id_right_identity.
  Qed.

  Lemma TrivialTriangle1_proper : forall X,
    (components_of (epsilon TrivialPreStable) (object_of (Susp TrivialPreStable) X) o 
     morphism_of (Susp TrivialPreStable) (components_of (eta TrivialPreStable) X))%morphism = 1%morphism.
  Proof.
    intro X.
    simpl.
    apply two_id_left_identity.
  Qed.

  Lemma TrivialTriangle2_proper : forall X,
    (morphism_of (Loop TrivialPreStable) (components_of (epsilon TrivialPreStable) X) o
     components_of (eta TrivialPreStable) (object_of (Loop TrivialPreStable) X))%morphism = 1%morphism.
  Proof.
    intro X.
    simpl.
    apply two_id_left_identity.
  Qed.

  Definition TrivialProperStable : ProperStableCategory.
  Proof.
    exact (Build_ProperStableCategory
      TrivialPreStable
      TrivialEta_is_iso_proper
      TrivialEpsilon_is_iso_proper
      TrivialTriangle1_proper
      TrivialTriangle2_proper).
  Defined.

  (** We have successfully constructed a trivial proper stable category.
      This example shows that the identity functor on any additive category
      can serve as both suspension and loop functors, yielding a proper stable
      structure where all the required isomorphisms are identities. *)

  End ChainComplexes.

  (** * Triangulated structure on TrivialProperStable *)

  Section TrivialTriangulated.
    Require Import Triangles PreStableCofiber.
    
    (** For any morphism in TwoCat, we need to define its cofiber *)
    Definition TrivialCofiber {X Y : SimpleBiproductCategory.TwoObj} 
      (f : morphism SimpleBiproductCategory.TwoCat X Y) : SimpleBiproductCategory.TwoObj.
    Proof.
      (* In our trivial category, the cofiber is always Zero *)
      exact SimpleBiproductCategory.Zero.
    Defined.

  (** The inclusion morphism from Y to cofiber(f) *)
    Definition TrivialCofiber_in {X Y : SimpleBiproductCategory.TwoObj} 
      (f : morphism SimpleBiproductCategory.TwoCat X Y) 
      : morphism SimpleBiproductCategory.TwoCat Y (TrivialCofiber f).
    Proof.
      unfold TrivialCofiber.
      destruct Y.
      - (* Y = Zero → Zero *)
        exact tt.
      - (* Y = One → Zero *)
        exact tt.
    Defined.

  (** The projection morphism from cofiber(f) to ΣX *)
    Definition TrivialCofiber_out {X Y : SimpleBiproductCategory.TwoObj} 
      (f : morphism SimpleBiproductCategory.TwoCat X Y) 
      : morphism SimpleBiproductCategory.TwoCat (TrivialCofiber f) (object_of TrivialSuspLoop X).
    Proof.
      unfold TrivialCofiber.
      simpl.
      (* Zero → X *)
      exact tt.
    Defined.

  (** Verify the first cofiber condition: cofiber_in ∘ f = 0 *)
    Lemma TrivialCofiber_cond1 {X Y : SimpleBiproductCategory.TwoObj} 
      (f : morphism SimpleBiproductCategory.TwoCat X Y) :
      (TrivialCofiber_in f o f)%morphism = 
      add_zero_morphism TwoCatAdditive.TwoAdditive X (TrivialCofiber f).
    Proof.
      unfold add_zero_morphism, zero_morphism.
      simpl.
      destruct X, Y; destruct f; reflexivity.
    Qed.

  (** Verify the second cofiber condition: cofiber_out ∘ cofiber_in = 0 *)
    Lemma TrivialCofiber_cond2 {X Y : SimpleBiproductCategory.TwoObj} 
      (f : morphism SimpleBiproductCategory.TwoCat X Y) :
      (TrivialCofiber_out f o TrivialCofiber_in f)%morphism = 
      add_zero_morphism TwoCatAdditive.TwoAdditive Y (object_of TrivialSuspLoop X).
    Proof.
      unfold add_zero_morphism, zero_morphism.
      simpl.
      destruct X, Y; destruct f; reflexivity.
    Qed.

  (** Verify the third cofiber condition: Σf ∘ cofiber_out = 0 *)
    Lemma TrivialCofiber_cond3 {X Y : SimpleBiproductCategory.TwoObj} 
      (f : morphism SimpleBiproductCategory.TwoCat X Y) :
      (morphism_of TrivialSuspLoop f o TrivialCofiber_out f)%morphism = 
      add_zero_morphism TwoCatAdditive.TwoAdditive (TrivialCofiber f) (object_of TrivialSuspLoop Y).
    Proof.
      unfold add_zero_morphism, zero_morphism.
      simpl.
      destruct X, Y; destruct f; reflexivity.
    Qed.

  (** Package the trivial cofiber structure *)
    Definition TrivialPreStableWithCofiber : PreStableCategoryWithCofiber.
    Proof.
      refine (Build_PreStableCategoryWithCofiber
        TrivialPreStable
        (fun X Y f => TrivialCofiber f)
        (fun X Y f => TrivialCofiber_in f)
        (fun X Y f => TrivialCofiber_out f)
        _ _ _).
      - (* cofiber_cond1 *)
        intros X Y f.
        apply TrivialCofiber_cond1.
      - (* cofiber_cond2 *)
        intros X Y f.
        apply TrivialCofiber_cond2.
      - (* cofiber_cond3 *)
        intros X Y f.
        apply TrivialCofiber_cond3.
    Defined.

  (** Every morphism extends to a distinguished triangle *)
    Lemma TrivialTR1 {X Y : SimpleBiproductCategory.TwoObj} 
      (f : morphism SimpleBiproductCategory.TwoCat X Y) :
      DistinguishedTriangle TrivialPreStable.
    Proof.
      apply (cofiber_triangle_distinguished TrivialPreStableWithCofiber f).
    Qed.

  (** Example: The distinguished triangle from the identity morphism *)
    Example identity_triangle : DistinguishedTriangle TrivialPreStable.
    Proof.
      apply (TrivialTR1 (1%morphism : morphism SimpleBiproductCategory.TwoCat 
                                       SimpleBiproductCategory.One 
                                       SimpleBiproductCategory.One)).
    Qed.

  (** Let's construct a concrete triangle example instead *)
    Definition concrete_triangle_example : Triangle TrivialPreStable.
    Proof.
      apply (@triangle_from_morphism TrivialPreStableWithCofiber
              SimpleBiproductCategory.One 
              SimpleBiproductCategory.One).
      exact 1%morphism.
    Defined.

  (** This concrete triangle is distinguished *)
    Lemma concrete_triangle_is_distinguished : 
      DistinguishedTriangle TrivialPreStable.
    Proof.
      apply (@cofiber_triangle_distinguished TrivialPreStableWithCofiber
              SimpleBiproductCategory.One 
              SimpleBiproductCategory.One).
      exact 1%morphism.
    Qed.

  Require Import TriangleRotation.

  (** Verify that rotation preserves distinguished triangles in our example *)
    Lemma concrete_triangle_rotation_distinguished : 
      DistinguishedTriangle TrivialPreStable.
    Proof.
      apply rotate_distinguished.
      apply concrete_triangle_is_distinguished.
    Qed.

  (** The trivial category satisfies the octahedral axiom trivially *)
    Lemma TrivialTR4_holds : 
      forall (X Y Z : object TrivialPreStable) 
             (f : morphism TrivialPreStable X Y) 
             (g : morphism TrivialPreStable Y Z),
      exists (u : morphism TrivialPreStable (TrivialCofiber f) (TrivialCofiber g)),
      (u o TrivialCofiber_in f)%morphism = (TrivialCofiber_in g o g)%morphism.
    Proof.
      intros X Y Z f g.
      (* In the trivial category, all cofibers are Zero *)
      exists tt.
      destruct X, Y, Z; destruct f; destruct g; reflexivity.
    Qed.

  (** We have shown that TrivialProperStable forms a triangulated category:
        - It has a cofiber structure (TrivialPreStableWithCofiber)
        - Every morphism extends to a distinguished triangle (TR1)
        - Distinguished triangles can be rotated (TR3)
        - The octahedral axiom holds (TR4)
        
        This is the simplest possible example where all functors are identity
        and all cofibers are the zero object. *)

  End TrivialTriangulated.

  (** * A non-trivial example: Graded abelian groups *)

  Section GradedAbelianGroups.
    Context `{Funext}.
    
    (** For simplicity, we'll use nat-graded groups *)
    Record GradedAbelianGroup := {
      graded_component : nat -> AbelianGroupWithLaws
    }.
    
    (** Morphisms are families of group homomorphisms *)
    Record GradedMorphism (G H : GradedAbelianGroup) := {
      graded_mor_component : forall (n : nat), 
        GroupHom (graded_component G n) (graded_component H n)
    }.

  (** Identity morphism *)
    Definition graded_id (G : GradedAbelianGroup) : GradedMorphism G G.
    Proof.
      refine (Build_GradedMorphism G G _).
      intro n.
      exact (id_hom (graded_component G n)).
    Defined.

  (** Composition of morphisms *)
    Definition graded_comp {A B C : GradedAbelianGroup} 
      (g : GradedMorphism B C) (f : GradedMorphism A B) : GradedMorphism A C.
    Proof.
      refine (Build_GradedMorphism A C _).
      intro n.
      exact (comp_hom (graded_mor_component B C g n) (graded_mor_component A B f n)).
    Defined.

  (** Morphisms are equal if their components are equal *)
    Lemma GradedMorphism_eq {G K : GradedAbelianGroup} (f g : GradedMorphism G K) :
      (forall n, graded_mor_component G K f n = graded_mor_component G K g n) -> f = g.
    Proof.
      intro Heq.
      destruct f as [f_comp].
      destruct g as [g_comp].
      simpl in Heq.
      f_ap.
      apply path_forall.
      exact Heq.
    Qed.

  (** The category of graded abelian groups *)
    Definition GradedAbGroupCat : PreCategory.
    Proof.
      refine (@Build_PreCategory
        GradedAbelianGroup
        GradedMorphism
        graded_id
        (@graded_comp)
        _ _ _ _).
      - (* associativity *)
        intros A B C D f g h.
        apply GradedMorphism_eq.
        intro n.
        simpl.
        symmetry.
        apply comp_hom_assoc.
      - (* left identity *)
        intros A B f.
        apply GradedMorphism_eq.
        intro n.
        simpl.
        apply comp_hom_id_left.
      - (* right identity *)
        intros A B f.
        apply GradedMorphism_eq.
        intro n.
        simpl.
        apply comp_hom_id_right.
      - (* truncation: morphisms form a set *)
        intros s d.
        apply (istrunc_equiv_istrunc _ 
          (equiv_adjointify
            (graded_mor_component s d)
            (Build_GradedMorphism s d)
            (fun f => idpath)
            (fun f => match f with Build_GradedMorphism comp => idpath end))^-1).
    Defined.

  (** The zero graded abelian group *)
    Definition ZeroGradedGroup : GradedAbelianGroup.
    Proof.
      refine (Build_GradedAbelianGroup _).
      intro n.
      exact TrivialGroup.
    Defined.

  (** ZeroGradedGroup is the zero object *)
    Theorem ZeroGradedGroup_is_zero : ZeroObject GradedAbGroupCat.
    Proof.
      refine (Build_ZeroObject GradedAbGroupCat ZeroGradedGroup _ _).
      - (* initial *)
        intro Y.
        apply Build_Contr with 
          (center := Build_GradedMorphism ZeroGradedGroup Y (fun n => zero_hom _ _)).
        intro f.
        apply GradedMorphism_eq.
        intro n.
        apply GroupHom_eq.
        apply path_forall. intro x.
        destruct x.
        simpl.
        symmetry.
        exact (hom_zero _ _ (graded_mor_component _ _ f n)).
      - (* terminal *)
        intro X.
        apply Build_Contr with
          (center := Build_GradedMorphism X ZeroGradedGroup (fun n => zero_hom _ _)).
        intro f.
        apply GradedMorphism_eq.
        intro n.
        apply GroupHom_eq.
        apply path_forall. intro x.
        destruct (hom_map _ _ (graded_mor_component _ _ f n) x).
        reflexivity.
    Defined.

  (** The shift functor on graded abelian groups *)
    Definition ShiftGradedGroup (G : GradedAbelianGroup) : GradedAbelianGroup.
    Proof.
      refine (Build_GradedAbelianGroup _).
      intro n.
      exact (graded_component G (S n)).
    Defined.

  (** The shift functor on morphisms *)
    Definition ShiftGradedMorphism {G K : GradedAbelianGroup} 
      (f : GradedMorphism G K) : GradedMorphism (ShiftGradedGroup G) (ShiftGradedGroup K).
    Proof.
      refine (Build_GradedMorphism _ _ _).
      intro n.
      exact (graded_mor_component G K f (S n)).
    Defined.

  (** Package shift as a functor *)
    Definition ShiftGradedFunctor : Functor GradedAbGroupCat GradedAbGroupCat.
    Proof.
      refine (Build_Functor 
        GradedAbGroupCat GradedAbGroupCat
        ShiftGradedGroup
        (@ShiftGradedMorphism)
        _ _).
      - (* composition *)
        intros G K L f g.
        apply GradedMorphism_eq.
        intro n.
        reflexivity.
      - (* identity *)
        intro G.
        apply GradedMorphism_eq.
        intro n.
        reflexivity.
    Defined.

Definition LoopGradedGroup (G : GradedAbelianGroup) : GradedAbelianGroup.
  Proof.
    refine (Build_GradedAbelianGroup _).
    intro n.
    destruct n as [|n'].
    - exact (graded_component G 0).
    - exact (graded_component G n').
  Defined.

Definition LoopGradedMorphism {G K : GradedAbelianGroup} 
    (f : GradedMorphism G K) : GradedMorphism (LoopGradedGroup G) (LoopGradedGroup K).
  Proof.
    refine (Build_GradedMorphism _ _ _).
    intro n.
    destruct n as [|n'].
    - exact (graded_mor_component G K f 0).
    - exact (graded_mor_component G K f n').
  Defined.

Definition LoopGradedFunctor : Functor GradedAbGroupCat GradedAbGroupCat.
  Proof.
    refine (Build_Functor 
      GradedAbGroupCat GradedAbGroupCat
      LoopGradedGroup
      (@LoopGradedMorphism)
      _ _).
    - intros G K L f g.
      apply GradedMorphism_eq.
      intro n.
      destruct n as [|n'].
      + reflexivity.
      + reflexivity.
    - intro G.
      apply GradedMorphism_eq.
      intro n.
      destruct n as [|n'].
      + reflexivity.
      + reflexivity.
  Defined.

Definition eta_graded_component (G : GradedAbelianGroup) 
    : GradedMorphism G (LoopGradedGroup (ShiftGradedGroup G)).
  Proof.
    refine (Build_GradedMorphism _ _ _).
    intro n.
    simpl.
    (* (Loop(Shift(G)))_n = match n with 0 => (Shift G)_0 = G_1 | S n' => (Shift G)_{n'} = G_{S n'} *)
    destruct n as [|n'].
    - (* degree 0: G_0 → G_1 - we need a morphism here *)
      exact (zero_hom (graded_component G 0) (graded_component G 1)).
    - (* degree S n': G_{S n'} → G_{S n'} *)
      exact (id_hom (graded_component G (S n'))).
  Defined.

Lemma eta_graded_natural {G K : GradedAbelianGroup} (f : GradedMorphism G K) :
    graded_comp (LoopGradedMorphism (ShiftGradedMorphism f)) (eta_graded_component G) =
    graded_comp (eta_graded_component K) f.
  Proof.
    apply GradedMorphism_eq.
    intro n.
    destruct n as [|n'].
    - (* degree 0 *)
      simpl.
      rewrite comp_zero_hom_left.
      rewrite comp_zero_hom_right.
      reflexivity.
    - (* degree S n' *)
      simpl.
      rewrite comp_hom_id_right.
      rewrite comp_hom_id_left.
      reflexivity.
  Qed.

Definition eta_graded : NaturalTransformation 
    (1%functor : Functor GradedAbGroupCat GradedAbGroupCat)
    ((LoopGradedFunctor o ShiftGradedFunctor)%functor).
  Proof.
    refine (Build_NaturalTransformation 
      (1%functor : Functor GradedAbGroupCat GradedAbGroupCat)
      ((LoopGradedFunctor o ShiftGradedFunctor)%functor)
      eta_graded_component _).
    intros G K f.
    simpl.
    symmetry.
    apply eta_graded_natural.
  Defined.

Definition epsilon_graded_component (G : GradedAbelianGroup) 
    : GradedMorphism (ShiftGradedGroup (LoopGradedGroup G)) G.
  Proof.
    refine (Build_GradedMorphism _ _ _).
    intro n.
    simpl.
    (* (Shift(Loop(G)))_n = (Loop(G))_{S n} *)
    (* When n = 0: (Loop G)_1 = G_0, so G_0 → G_0 *)
    (* When n = S n': (Loop G)_{S (S n')} = G_{S n'}, so G_{S n'} → G_{S n'} *)
    exact (id_hom _).
  Defined.

Lemma epsilon_graded_natural {G K : GradedAbelianGroup} (f : GradedMorphism G K) :
    graded_comp f (epsilon_graded_component G) =
    graded_comp (epsilon_graded_component K) (ShiftGradedMorphism (LoopGradedMorphism f)).
  Proof.
    apply GradedMorphism_eq.
    intro n.
    simpl.
    rewrite comp_hom_id_left.
    rewrite comp_hom_id_right.
    reflexivity.
  Qed.

Definition epsilon_graded : NaturalTransformation 
    ((ShiftGradedFunctor o LoopGradedFunctor)%functor)
    (1%functor : Functor GradedAbGroupCat GradedAbGroupCat).
  Proof.
    refine (Build_NaturalTransformation 
      ((ShiftGradedFunctor o LoopGradedFunctor)%functor)
      (1%functor : Functor GradedAbGroupCat GradedAbGroupCat)
      epsilon_graded_component _).
    intros G K f.
    simpl.
    symmetry.
    apply epsilon_graded_natural.
  Defined.

Definition DirectSumGraded (G K : GradedAbelianGroup) : GradedAbelianGroup.
  Proof.
    refine (Build_GradedAbelianGroup _).
    intro n.
    exact (DirectSum (graded_component G n) (graded_component K n)).
  Defined.


Lemma loop_graded_preserves_biproduct (G K : GradedAbelianGroup) :
    LoopGradedGroup (DirectSumGraded G K) = 
    DirectSumGraded (LoopGradedGroup G) (LoopGradedGroup K).
  Proof.
    unfold LoopGradedGroup, DirectSumGraded.
    f_ap.
    apply path_forall. intro n.
    destruct n as [|n'].
    - reflexivity.
    - reflexivity.
  Qed.

Definition graded_inj1 (G K : GradedAbelianGroup) : GradedMorphism G (DirectSumGraded G K).
  Proof.
    refine (Build_GradedMorphism _ _ _).
    intro n.
    exact (inj1 (graded_component G n) (graded_component K n)).
  Defined.

  Definition graded_inj2 (G K : GradedAbelianGroup) : GradedMorphism K (DirectSumGraded G K).
  Proof.
    refine (Build_GradedMorphism _ _ _).
    intro n.
    exact (inj2 (graded_component G n) (graded_component K n)).
  Defined.

  Definition graded_proj1 (G K : GradedAbelianGroup) : GradedMorphism (DirectSumGraded G K) G.
  Proof.
    refine (Build_GradedMorphism _ _ _).
    intro n.
    exact (proj1 (graded_component G n) (graded_component K n)).
  Defined.

  Definition graded_proj2 (G K : GradedAbelianGroup) : GradedMorphism (DirectSumGraded G K) K.
  Proof.
    refine (Build_GradedMorphism _ _ _).
    intro n.
    exact (proj2 (graded_component G n) (graded_component K n)).
  Defined.

  Lemma graded_beta_l (G K : GradedAbelianGroup) : 
    graded_comp (graded_proj1 G K) (graded_inj1 G K) = graded_id G.
  Proof.
    apply GradedMorphism_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro x.
    reflexivity.
  Qed.

  Lemma graded_beta_r (G K : GradedAbelianGroup) : 
    graded_comp (graded_proj2 G K) (graded_inj2 G K) = graded_id K.
  Proof.
    apply GradedMorphism_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro x.
    reflexivity.
  Qed.

  Lemma graded_mixed_l (G K : GradedAbelianGroup) : 
    graded_comp (graded_proj1 G K) (graded_inj2 G K) = 
    Build_GradedMorphism K G (fun n => zero_hom _ _).
  Proof.
    apply GradedMorphism_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro x.
    reflexivity.
  Qed.

Lemma graded_mixed_r (G K : GradedAbelianGroup) : 
    graded_comp (graded_proj2 G K) (graded_inj1 G K) = 
    Build_GradedMorphism G K (fun n => zero_hom _ _).
  Proof.
    apply GradedMorphism_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro x.
    reflexivity.
  Qed.

  Definition graded_coprod_mor (G K W : GradedAbelianGroup) 
    (f : GradedMorphism G W) (g : GradedMorphism K W) 
    : GradedMorphism (DirectSumGraded G K) W.
  Proof.
    refine (Build_GradedMorphism _ _ _).
    intro n.
    set (fn := graded_mor_component G W f n).
    set (gn := graded_mor_component K W g n).
    refine (Build_GroupHom (DirectSum (graded_component G n) (graded_component K n))
                          (graded_component W n)
                          (fun p => plus (group (graded_component W n))
                                        (hom_map _ _ fn (fst p))
                                        (hom_map _ _ gn (snd p))) _ _).
    - simpl.
      rewrite (hom_zero _ _ fn).
      rewrite (hom_zero _ _ gn).
      apply (plus_zero_l _ (laws (graded_component W n))).
    - intros p1 p2.
      simpl.
      rewrite (hom_plus _ _ fn).
      rewrite (hom_plus _ _ gn).
      set (fx1 := hom_map _ _ fn (fst p1)).
      set (fx2 := hom_map _ _ fn (fst p2)).
      set (gy1 := hom_map _ _ gn (snd p1)).
      set (gy2 := hom_map _ _ gn (snd p2)).
      rewrite <- (plus_assoc _ (laws (graded_component W n)) fx1 gy1 _).
      rewrite (plus_assoc _ (laws (graded_component W n)) gy1 fx2 gy2).
      rewrite (plus_comm _ (laws (graded_component W n)) gy1 fx2).
      rewrite <- (plus_assoc _ (laws (graded_component W n)) fx2 gy1 gy2).
      rewrite (plus_assoc _ (laws (graded_component W n)) fx1 fx2 _).
      reflexivity.
  Defined.

Lemma graded_coprod_beta_l (G K W : GradedAbelianGroup) 
    (f : GradedMorphism G W) (g : GradedMorphism K W) :
    graded_comp (graded_coprod_mor G K W f g) (graded_inj1 G K) = f.
  Proof.
    apply GradedMorphism_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro x.
    simpl.
    rewrite (hom_zero _ _ (graded_mor_component K W g n)).
    apply (plus_zero_r _ (laws (graded_component W n))).
  Qed.

  Lemma graded_coprod_beta_r (G K W : GradedAbelianGroup) 
    (f : GradedMorphism G W) (g : GradedMorphism K W) :
    graded_comp (graded_coprod_mor G K W f g) (graded_inj2 G K) = g.
  Proof.
    apply GradedMorphism_eq.
    intro n.
    simpl.
    apply GroupHom_eq.
    apply path_forall. intro x.
    simpl.
    rewrite (hom_zero _ _ (graded_mor_component G W f n)).
    apply (plus_zero_l _ (laws (graded_component W n))).
  Qed.

  Definition graded_prod_mor (W G K : GradedAbelianGroup) 
    (f : GradedMorphism W G) (g : GradedMorphism W K) 
    : GradedMorphism W (DirectSumGraded G K).
  Proof.
    refine (Build_GradedMorphism _ _ _).
    intro n.
    refine (Build_GroupHom (graded_component W n)
                          (DirectSum (graded_component G n) (graded_component K n))
                          (fun w => (hom_map _ _ (graded_mor_component W G f n) w,
                                    hom_map _ _ (graded_mor_component W K g n) w)) _ _).
    - simpl.
      f_ap.
      * apply (hom_zero _ _ (graded_mor_component W G f n)).
      * apply (hom_zero _ _ (graded_mor_component W K g n)).
    - intros w1 w2.
      simpl.
      f_ap.
      * apply (hom_plus _ _ (graded_mor_component W G f n)).
      * apply (hom_plus _ _ (graded_mor_component W K g n)).
  Defined.

  Lemma graded_prod_beta_l (W G K : GradedAbelianGroup) 
    (f : GradedMorphism W G) (g : GradedMorphism W K) :
    graded_comp (graded_proj1 G K) (graded_prod_mor W G K f g) = f.
  Proof.
    apply GradedMorphism_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intro w.
    reflexivity.
  Qed.

 Lemma graded_prod_beta_r (W G K : GradedAbelianGroup) 
    (f : GradedMorphism W G) (g : GradedMorphism W K) :
    graded_comp (graded_proj2 G K) (graded_prod_mor W G K f g) = g.
  Proof.
    apply GradedMorphism_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intro w.
    reflexivity.
  Qed.

  Lemma graded_zero_morphism_eq (G K : GradedAbelianGroup) :
    zero_morphism ZeroGradedGroup_is_zero G K = 
    Build_GradedMorphism G K (fun n => zero_hom _ _).
  Proof.
    unfold zero_morphism.
    simpl.
    apply GradedMorphism_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intro x.
    reflexivity.
  Qed.

  Global Instance GradedMorphism_IsHSet `{Funext} (G K : GradedAbelianGroup) 
    : IsHSet (GradedMorphism G K).
  Proof.
    assert (equiv_to_prod : GradedMorphism G K <~> 
      forall n, GroupHom (graded_component G n) (graded_component K n)).
    {
      apply (equiv_adjointify
        (graded_mor_component G K)
        (Build_GradedMorphism G K)).
      - intro f.
        apply path_forall. intro n.
        reflexivity.
      - intros [comp].
        reflexivity.
    }
    apply (istrunc_equiv_istrunc _ equiv_to_prod^-1).
  Qed.

  Lemma graded_coprod_unique (G K W : GradedAbelianGroup) 
    (f : GradedMorphism G W) (g : GradedMorphism K W)
    (h : GradedMorphism (DirectSumGraded G K) W) :
    graded_comp h (graded_inj1 G K) = f ->
    graded_comp h (graded_inj2 G K) = g ->
    h = graded_coprod_mor G K W f g.
  Proof.
    intros Hl Hr.
    apply GradedMorphism_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intros [x y].
    assert (Hxy_decomp : (x, y) = 
      plus (group (DirectSum (graded_component G n) (graded_component K n)))
           (x, zero (group (graded_component K n)))
           (zero (group (graded_component G n)), y)).
    {
      simpl.
      f_ap.
      - symmetry. apply (plus_zero_r _ (laws (graded_component G n))).
      - symmetry. apply (plus_zero_l _ (laws (graded_component K n))).
    }
    rewrite Hxy_decomp.
    rewrite (hom_plus _ _ (graded_mor_component _ _ h n)).
    pose proof (ap (fun k => graded_mor_component _ _ k n) Hl) as Hl_n.
    pose proof (ap (fun k => graded_mor_component _ _ k n) Hr) as Hr_n.
    simpl in *.
    assert (Hlx : hom_map _ _ (graded_mor_component _ _ h n) 
                          (x, zero (group (graded_component K n))) =
                  hom_map _ _ (graded_mor_component G W f n) x).
    {
      change (hom_map _ _ (graded_mor_component _ _ h n) 
                     (hom_map _ _ (inj1 _ _) x) =
              hom_map _ _ (graded_mor_component G W f n) x).
      unfold comp_hom in Hl_n.
      exact (ap (fun k => hom_map _ _ k x) Hl_n).
    }
    assert (Hry : hom_map _ _ (graded_mor_component _ _ h n) 
                          (zero (group (graded_component G n)), y) =
                  hom_map _ _ (graded_mor_component K W g n) y).
    {
      change (hom_map _ _ (graded_mor_component _ _ h n) 
                     (hom_map _ _ (inj2 _ _) y) =
              hom_map _ _ (graded_mor_component K W g n) y).
      unfold comp_hom in Hr_n.
      exact (ap (fun k => hom_map _ _ k y) Hr_n).
    }
    rewrite Hlx, Hry.
    simpl.
    f_ap.
    - rewrite (plus_zero_r _ (laws (graded_component G n))).
      reflexivity.
    - rewrite (plus_zero_l _ (laws (graded_component K n))).
      reflexivity.
  Qed.

  Lemma graded_prod_unique (W G K : GradedAbelianGroup) 
    (f : GradedMorphism W G) (g : GradedMorphism W K)
    (h : GradedMorphism W (DirectSumGraded G K)) :
    graded_comp (graded_proj1 G K) h = f ->
    graded_comp (graded_proj2 G K) h = g ->
    h = graded_prod_mor W G K f g.
  Proof.
    intros Hl Hr.
    apply GradedMorphism_eq.
    intro n.
    apply GroupHom_eq.
    apply path_forall. intro w.
    pose proof (ap (fun k => graded_mor_component _ _ k n) Hl) as Hl_n.
    pose proof (ap (fun k => graded_mor_component _ _ k n) Hr) as Hr_n.
    simpl in *.
    pose proof (ap (fun k => hom_map _ _ k w) Hl_n) as Hlw.
    pose proof (ap (fun k => hom_map _ _ k w) Hr_n) as Hrw.
    simpl in *.
    destruct (hom_map _ _ (graded_mor_component _ _ h n) w) as [a b].
    simpl in *.
    f_ap; assumption.
  Qed.

  Definition GradedBiproduct (G K : GradedAbelianGroup) 
    : @Biproduct GradedAbGroupCat G K ZeroGradedGroup_is_zero.
  Proof.
    pose (bdata := Build_BiproductData GradedAbGroupCat G K 
      (DirectSumGraded G K)
      (graded_inj1 G K)
      (graded_inj2 G K)
      (graded_proj1 G K)
      (graded_proj2 G K)).
    assert (bis : IsBiproduct bdata ZeroGradedGroup_is_zero).
    {
      simple refine (Build_IsBiproduct _ _ _ _ _ _ _ _ _).
      - apply graded_beta_l.
      - apply graded_beta_r.
      - simpl. rewrite graded_mixed_l. symmetry. apply graded_zero_morphism_eq.
      - simpl. rewrite graded_mixed_r. symmetry. apply graded_zero_morphism_eq.
    }
    assert (buni : HasBiproductUniversal bdata).
    {
      simple refine (Build_HasBiproductUniversal _ _ _ _ _ _).
      - intros W f g.
        apply (Build_Contr _ (graded_coprod_mor G K W f g; 
                             (graded_coprod_beta_l G K W f g, 
                              graded_coprod_beta_r G K W f g))).
        intros [h [Hl Hr]].
        apply path_sigma_uncurried.
        simpl.
        exists ((graded_coprod_unique G K W f g h Hl Hr)^).
        apply path_ishprop.
      - intros W f g.
        apply (Build_Contr _ (graded_prod_mor W G K f g; 
                             (graded_prod_beta_l W G K f g, 
                              graded_prod_beta_r W G K f g))).
        intros [h [Hl Hr]].
        apply path_sigma_uncurried.
        simpl.
        exists ((graded_prod_unique W G K f g h Hl Hr)^).
        apply path_ishprop.
    }
    exact (Build_Biproduct _ _ _ _ bdata bis buni).
  Defined.

  Definition GradedAdditive `{Funext} : AdditiveCategory.
  Proof.
    exact (Build_AdditiveCategory 
      GradedAbGroupCat
      ZeroGradedGroup_is_zero
      GradedBiproduct).
  Defined.

Lemma loop_graded_preserves_zero : 
    LoopGradedGroup ZeroGradedGroup = ZeroGradedGroup.
  Proof.
    unfold LoopGradedGroup, ZeroGradedGroup.
    f_ap.
    apply path_forall. intro n.
    destruct n; reflexivity.
  Qed.

Definition LoopGradedAdditiveFunctor `{Funext} : AdditiveFunctor GradedAdditive GradedAdditive.
  Proof.
    refine (Build_AdditiveFunctor 
      GradedAdditive GradedAdditive
      LoopGradedFunctor
      _ _).
    - (* preserves_zero *)
      exact loop_graded_preserves_zero.
    - (* preserves_biproduct *)
      exact loop_graded_preserves_biproduct.
  Defined.

Lemma shift_graded_preserves_zero : 
    ShiftGradedGroup ZeroGradedGroup = ZeroGradedGroup.
  Proof.
    unfold ShiftGradedGroup, ZeroGradedGroup.
    f_ap.
  Qed.

Lemma shift_graded_preserves_biproduct (G K : GradedAbelianGroup) :
    ShiftGradedGroup (DirectSumGraded G K) = 
    DirectSumGraded (ShiftGradedGroup G) (ShiftGradedGroup K).
  Proof.
    unfold ShiftGradedGroup, DirectSumGraded.
    f_ap.
  Qed.

Definition ShiftGradedAdditiveFunctor `{Funext} : AdditiveFunctor GradedAdditive GradedAdditive.
  Proof.
    refine (Build_AdditiveFunctor 
      GradedAdditive GradedAdditive
      ShiftGradedFunctor
      _ _).
    - (* preserves_zero *)
      exact shift_graded_preserves_zero.
    - (* preserves_biproduct *)
      exact shift_graded_preserves_biproduct.
  Defined.

Definition GradedPreStable `{Funext} : PreStableCategory.
  Proof.
    exact (Build_PreStableCategory
      GradedAdditive
      ShiftGradedAdditiveFunctor
      LoopGradedAdditiveFunctor
      eta_graded
      epsilon_graded).
  Defined.

Lemma graded_triangle_1 : forall G,
    graded_comp (epsilon_graded_component (ShiftGradedGroup G)) 
                (ShiftGradedMorphism (eta_graded_component G)) = 
    graded_id (ShiftGradedGroup G).
  Proof.
    intro G.
    apply GradedMorphism_eq.
    intro n.
    simpl.
    destruct n as [|n'].
    - (* degree 0: id ∘ id = id *)
      rewrite comp_hom_id_left.
      reflexivity.
    - (* degree S n': id ∘ id = id *)
      rewrite comp_hom_id_left.
      reflexivity.
  Qed.

Theorem graded_is_prestable `{Funext} : PreStableCategory.
  Proof.
    exact GradedPreStable.
  Qed.

Theorem shift_loop_compose_id `{Funext} (G : GradedAbelianGroup) :
    ShiftGradedGroup (LoopGradedGroup G) = G.
  Proof.
    unfold ShiftGradedGroup, LoopGradedGroup.
    destruct G as [g].
    simpl.
    f_ap.
  Qed.
