(** * Wedge Sums Preserve Connectivity in HoTT
    
    This module proves that wedge sums (coproducts in the category of pointed 
    types) preserve n-connectedness. This fundamental result appears to be 
    original in the context of synthetic homotopy theory.
    
    Author: Charles Norton
    Date: July 6th 2025
    License: GNU Lesser General Public License Version 2.1
    
    Compatibility: HoTT library (Coq 8.16+)
*)

Require Import HoTT.Basics.
Require Import HoTT.Types.
Require Import HoTT.Pointed.Core.
Require Import HoTT.Truncations.Core.
Require Import HoTT.Truncations.Connectedness.
Require Import HoTT.Colimits.Pushout.

(** ** Overview
    
    The wedge sum X ∨ Y of two pointed types is their coproduct in the category
    of pointed types. It is constructed by taking the disjoint union and 
    identifying the basepoints.
    
    A type is n-connected if its n-truncation is contractible. This module 
    establishes that if X and Y are n-connected pointed types, then their 
    wedge sum X ∨ Y is also n-connected.
    
    While this is a standard result in classical homotopy theory, formalizing 
    it synthetically in HoTT requires careful management of:
    
    - Higher inductive types (pushouts)
    - Truncation levels and connectivity
    - Path algebra and coherence conditions
    - The interplay between pointed types and their underlying types
    
    This formalization provides a foundation for more advanced results in 
    synthetic homotopy theory that use wedge constructions.
*)

(** ** Construction of Wedge Sums
    
    We construct the wedge sum as a pushout (a special case of a coequalizer).
    Given pointed types (X, x₀) and (Y, y₀), we form the pushout of the 
    diagram:
    
        unit_name x₀ : Unit → X
        unit_name y₀ : Unit → Y
    
    This identifies x₀ and y₀ in the disjoint union X + Y.
*)

(** Helper functions that constantly return the basepoints *)
Definition wedge_f (X Y : pType) : Unit -> X := fun _ => point X.
Definition wedge_g (X Y : pType) : Unit -> Y := fun _ => point Y.

(** The carrier type of a wedge sum as a pushout *)
Definition Wedge (X Y : pType) : Type :=
  Pushout (unit_name (point X)) (unit_name (point Y)).

(** The wedge sum as a pointed type, with basepoint from the left injection *)
Definition pWedge (X Y : pType) : pType :=
  Build_pType (Wedge X Y) (pushl (point X)).

(** ** Basic Properties of Wedge Sums *)

(** The basepoint of the wedge is the left injection of X's basepoint *)
Lemma wedge_point (X Y : pType) : point (pWedge X Y) = pushl (point X).
Proof.
  reflexivity.
Qed.

(** The glue path identifies the two basepoints *)
Lemma wedge_glue (X Y : pType) : 
  pushl (point X) = pushr (point Y) :> Wedge X Y.
Proof.
  exact (pglue tt).
Qed.

(** Alternative name for the glue path *)
Lemma wedge_glue_basepoints (X Y : pType) :
  pushl (point X) = pushr (point Y) :> Wedge X Y.
Proof.
  exact (pglue tt).
Qed.

(** ** Elimination Principle for Wedges
    
    To define a function out of a wedge, we need:
    - A function on X
    - A function on Y  
    - A proof that they agree on the basepoints (up to transport)
*)
Definition wedge_ind {X Y : pType} (P : Wedge X Y -> Type)
  (f : forall x : X, P (pushl x))
  (g : forall y : Y, P (pushr y))
  (p : transport P (pglue tt) (f (point X)) = g (point Y)) :
  forall w : Wedge X Y, P w.
Proof.
  refine (Pushout_ind P f g _).
  intro u; destruct u.
  exact p.
Defined.

(** ** Technical Lemmas about Unit and Basepoints
    
    Since our pushout uses unit_name to make Unit → X functions,
    we need several lemmas about how unit_name behaves.
*)

(** unit_name always returns the same point regardless of input *)
Lemma unit_name_constant {A : Type} (a : A) (u u' : Unit) :
  unit_name a u = unit_name a u'.
Proof.
  destruct u, u'. reflexivity.
Qed.

(** Left injection of unit_name gives the basepoint *)
Lemma pushl_unit_name_point (X Y : pType) (u : Unit) :
  pushl (unit_name (point X) u) = pushl (point X) :> Wedge X Y.
Proof.
  destruct u. reflexivity.
Qed.

(** Alternative formulation *)
Lemma pushl_unit_name_eq (X Y : pType) (u : Unit) :
  pushl (unit_name (point X) u) = pushl (point X) :> Wedge X Y.
Proof.
  destruct u. reflexivity.
Qed.

(** Right injection of unit_name gives the basepoint *)
Lemma pushr_unit_name_point (X Y : pType) (u : Unit) :
  pushr (unit_name (point Y) u) = pushr (point Y) :> Wedge X Y.
Proof.
  destruct u. reflexivity.
Qed.

(** All left elements from Unit map to the same point *)
Lemma wedge_pushl_all_equal (X Y : pType) (u : Unit) :
  pushl (unit_name (point X) u) = pushl (point X) :> Wedge X Y.
Proof.
  destruct u. reflexivity.
Qed.

(** All right elements from Unit map to the same point *)
Lemma wedge_pushr_all_equal (X Y : pType) (u : Unit) :
  pushr (unit_name (point Y) u) = pushr (point Y) :> Wedge X Y.
Proof.
  destruct u. reflexivity.
Qed.

(** The pglue path for any unit element *)
Lemma wedge_pglue_eq (X Y : pType) (u : Unit) :
  pushl (point X) = pushr (point Y) :> Wedge X Y.
Proof.
  exact (pglue u).
Qed.

(** ** Truncation and Connectivity Lemmas *)

(** Truncation preserves paths *)
Lemma tr_path {n : trunc_index} {A : Type} {x y : A} (p : x = y) :
  tr x = tr y :> Tr n A.
Proof.
  exact (ap tr p).
Qed.

(** In an n-connected type, all truncated elements are equal *)
Lemma tr_eq_of_connected {n : trunc_index} {A : Type} 
  (HA : IsConnected n A) (a b : A) :
  tr a = tr b :> Tr n A.
Proof.
  apply path_contr.
Qed.

(** Special case for 0-connected types *)
Lemma connected_implies_tr_equal {A : Type} 
  (HA : IsConnected 0 A) (a b : A) :
  tr a = tr b :> Tr 0 A.
Proof.
  apply path_contr.
Qed.

(** ** Transport Lemmas for Path Types
    
    These lemmas help manage transport in path types, which appears
    frequently when working with pushout induction.
*)

(** Transport in a pushout *)
Lemma transport_paths_pushout_pglue {A B C : Type} {f : B -> A} {g : B -> C} 
  (P : Pushout f g -> Type) (Q : forall w, P w) (b : B) :
  transport P (pglue b) (Q (pushl (f b))) = Q (pushr (g b)).
Proof.
  apply apD.
Qed.

(** Transport for paths with constant right-hand side *)
Lemma transport_paths_r_constant {A : Type} {n : trunc_index} 
  {x1 x2 : A} (p : x1 = x2) (y : Tr n A) (q : tr x1 = y) :
  transport (fun x => tr x = y) p q = ap tr p^ @ q.
Proof.
  destruct p. simpl. 
  rewrite concat_1p.
  reflexivity.
Qed.

(** Specific transport computation for our wedge case *)
Lemma transport_wedge_truncation_eq (n : trunc_index) (X Y : pType) :
  transport (fun w : Wedge X Y => tr w = tr (pushl (point X)) :> Tr n (Wedge X Y)) 
    (pglue tt)
    (1 : tr (pushl (point X)) = tr (pushl (point X)))
  = ap tr (pglue tt)^.
Proof.
  rewrite transport_paths_FlFr.
  rewrite ap_V.
  rewrite concat_p1.
  assert (H : ap (fun _ : Wedge X Y => tr (pushl (point X)) : Tr n (Wedge X Y)) (pglue tt) = 1).
  { apply ap_const. }
  rewrite H.
  exact (concat_p1 _).
Qed.

(** ** Main Connectivity Preservation Proof
    
    The proof strategy:
    1. Show that the n-truncation of the wedge has a center: tr(pushl(point X))
    2. Show that every truncated element equals this center
    3. Use pushout induction to handle left, right, and glue cases
    4. Carefully manage the coherence condition
*)

(** The center of the wedge truncation *)
Definition wedge_truncation_center (n : trunc_index) (X Y : pType) : Tr n (Wedge X Y) :=
  tr (point (pWedge X Y)).

(** The truncation of the basepoint equals the center *)
Lemma wedge_truncation_basepoint (n : trunc_index) (X Y : pType) :
  wedge_truncation_center n X Y = tr (pushl (point X)) :> Tr n (Wedge X Y).
Proof.
  reflexivity.
Qed.

(** For the pushout from Unit, left elements give reflexivity *)
Definition wedge_left_case (n : trunc_index) (X Y : pType) (x : Unit) :
  tr (pushl (unit_name (point X) x)) = tr (pushl (point X)) :> Tr n (Wedge X Y).
Proof.
  destruct x. reflexivity.
Defined.

(** For the pushout from Unit, right elements connect via the glue *)
Definition wedge_right_case (n : trunc_index) (X Y : pType) (y : Unit) :
  tr (pushr (unit_name (point Y) y)) = tr (pushl (point X)) :> Tr n (Wedge X Y).
Proof.
  destruct y. exact (ap tr (pglue tt)^).
Defined.

(** The coherence condition: left and right cases agree on the glue *)
Lemma wedge_glue_coherence (n : trunc_index) (X Y : pType) (u : Unit) :
  transport (fun w : Wedge X Y => tr w = tr (pushl (point X)) :> Tr n (Wedge X Y))
    (pglue u)
    (wedge_left_case n X Y u) = 
  wedge_right_case n X Y u.
Proof.
  destruct u.
  unfold wedge_left_case, wedge_right_case.
  simpl.
  exact (transport_wedge_truncation_eq n X Y).
Qed.

(** ** Connectivity Lemmas for Components
    
    These lemmas show that if X (or Y) is n-connected, then all elements
    from X (or Y) have equal truncations in the wedge.
*)

(** For n-connected X, all left elements have equal truncations *)
Lemma tr_pushl_connected {n : trunc_index} {X Y : pType} 
  (HX : IsConnected n X) (x : X) :
  tr (pushl x) = tr (pushl (point X)) :> Tr n (Wedge X Y).
Proof.
  (* Use functoriality of truncation *)
  exact (ap (Trunc_functor n pushl) (path_contr (tr x) (tr (point X)))).
Defined.

(** For n-connected Y, all right elements have equal truncations *)
Lemma tr_pushr_connected {n : trunc_index} {X Y : pType} 
  (HY : IsConnected n Y) (y : Y) :
  tr (pushr y) = tr (pushl (point X)) :> Tr n (Wedge X Y).
Proof.
  (* First show tr (pushr y) = tr (pushr (point Y)) *)
  transitivity (tr (pushr (point Y)) : Tr n (Wedge X Y)).
  - exact (ap (Trunc_functor n (@pushr _ _ _ (unit_name (point X)) (unit_name (point Y)))) 
              (path_contr (tr y) (tr (point Y)))).
  (* Then use the glue path *)
  - exact (ap tr (pglue tt)^).
Defined.

(** At the basepoint, tr_pushl_connected gives reflexivity *)
Lemma tr_pushl_connected_point (n : trunc_index) (X Y : pType) 
  (HX : IsConnected n X) :
  tr_pushl_connected (Y:=Y) HX (point X) = 1.
Proof.
  unfold tr_pushl_connected.
  (* In a contractible type, the canonical path to the center is 1 when start = end *)
  assert (H : @path_contr (Tr n X) HX (tr (point X)) (tr (point X)) = idpath _).
  { apply path_ishprop. }
  rewrite H.
  (* ap f 1 = 1 *)
  exact (ap_1 _ _).
Qed.

(** At the basepoint, tr_pushr_connected gives the glue path *)
Lemma tr_pushr_connected_point (n : trunc_index) (X Y : pType) 
  (HY : IsConnected n Y) :
  tr_pushr_connected (X:=X) HY (point Y) = ap tr (pglue tt)^.
Proof.
  unfold tr_pushr_connected.
  (* The first part: path_contr at the same point is 1 *)
  assert (H : @path_contr (Tr n Y) HY (tr (point Y)) (tr (point Y)) = idpath _).
  { apply path_ishprop. }
  rewrite H.
  rewrite (ap_1 _ _).
  (* 1 @ p = p *)
  apply concat_1p.
Qed.

(** The main coherence lemma for wedge truncation *)
Lemma wedge_truncation_coherence (n : trunc_index) (X Y : pType) 
  (HX : IsConnected n X) (HY : IsConnected n Y) (u : Unit) :
  transport (fun w => tr w = tr (pushl (point X)) :> Tr n (Wedge X Y))
    (pglue u)
    (tr_pushl_connected HX (unit_name (point X) u))
  = tr_pushr_connected HY (unit_name (point Y) u).
Proof.
  destruct u.
  (* Let's understand what transport does here *)
  rewrite transport_paths_FlFr.
  (* ap of constant function is 1 *)
  rewrite ap_const.
  (* Now simplify the concatenation with 1 *)
  rewrite concat_p1.
  (* Use our lemmas about the values at basepoints *)
  rewrite tr_pushl_connected_point.
  rewrite tr_pushr_connected_point.
  (* (ap tr (pglue tt))^ @ 1 = ap tr (pglue tt)^ *)
  rewrite concat_p1.
  (* We need to show (ap tr (pglue tt))^ = ap tr (pglue tt)^ *)
  rewrite ap_V.
  reflexivity.
Qed.

(** Any element of the wedge has its truncation equal to the center *)
Lemma wedge_truncation_eq_center (n : trunc_index) (X Y : pType) 
  (HX : IsConnected n X) (HY : IsConnected n Y) 
  (w : Wedge X Y) :
  tr w = tr (pushl (point X)) :> Tr n (Wedge X Y).
Proof.
  unfold Wedge in *.
  refine (Pushout_ind 
    (fun w => tr w = tr (pushl (point X)) :> Tr n _)
    (tr_pushl_connected HX)
    (tr_pushr_connected HY)
    _ w).
  - (* Coherence *)
    exact (wedge_truncation_coherence n X Y HX HY).
Defined.

(** ** Main Theorem
    
    The wedge sum of two n-connected pointed types is n-connected.
    
    This is proven by showing that the n-truncation of X ∨ Y is contractible,
    with center tr(pushl(point X)) and contraction given by 
    wedge_truncation_eq_center.
*)
Theorem wedge_preserves_connectedness (n : trunc_index) (X Y : pType)
  (HX : IsConnected n X) (HY : IsConnected n Y) :
  IsConnected n (pWedge X Y).
Proof.
  (* To show n-connectedness, we need to show Tr n (Wedge X Y) is contractible *)
  apply (Build_Contr _ (tr (pushl (point X)))).
  (* Every element equals the center *)
  intro x.
  strip_truncations.
  symmetry.
  apply wedge_truncation_eq_center.
  - exact HX.
  - exact HY.
Defined.

(** ** Examples and Applications *)

Require Import HoTT.Spaces.Circle.

(** *** Connectivity of the Circle
    
    We first establish that the circle is 0-connected, which will be used
    in several examples.
*)
Lemma circle_0_connected : IsConnected 0 Circle.
Proof.
  (* A type is 0-connected if its 0-truncation is contractible *)
  (* For the circle, we can show any two points are merely equal *)
  apply (Build_Contr _ (tr base)).
  intro x.
  strip_truncations.
  (* Use circle induction *)
  apply (Circle_ind (fun c => tr base = tr c) (idpath _)).
  (* Loop case: Need to show transport preserves the path *)
  apply path_ishprop.
Defined.

(** *** Example 1: Wedge of two circles
    
    The wedge S¹ ∨ S¹ (figure-eight) is 0-connected.
*)
Example wedge_circles_connected : 
  IsConnected 0 (pWedge (Build_pType Circle base) (Build_pType Circle base)).
Proof.
  apply wedge_preserves_connectedness.
  - exact circle_0_connected.
  - exact circle_0_connected.
Defined.

(** *** Example 2: Wedge with contractible type
    
    Wedging with a contractible type preserves connectivity.
*)
Example wedge_circle_unit_connected : 
  IsConnected 0 (pWedge (Build_pType Circle base) (Build_pType Unit tt)).
Proof.
  apply wedge_preserves_connectedness.
  - exact circle_0_connected.
  - (* Unit is 0-connected (actually contractible) *)
    apply contr_inhabited_hprop.
    + exact _.
    + apply tr. exact tt.
Defined.

(** *** Example 3: Triple wedge
    
    Connectivity is preserved under iterated wedging.
*)
Example wedge_three_circles_connected : 
  IsConnected 0 (pWedge (Build_pType Circle base) 
                        (pWedge (Build_pType Circle base) 
                                (Build_pType Circle base))).
Proof.
  apply wedge_preserves_connectedness.
  - exact circle_0_connected.
  - apply wedge_preserves_connectedness.
    + exact circle_0_connected.
    + exact circle_0_connected.
Defined.

(** *** Example 4: Bouquet of circles
    
    A bouquet of n circles is 0-connected for any n.
*)
Fixpoint bouquet_circles (n : nat) : pType :=
  match n with
  | O => Build_pType Unit tt
  | S n' => pWedge (Build_pType Circle base) (bouquet_circles n')
  end.

Lemma bouquet_circles_connected (n : nat) : IsConnected 0 (bouquet_circles n).
Proof.
  induction n.
  - (* Base case: Unit is 0-connected *)
    simpl.
    apply contr_inhabited_hprop.
    + exact _.
    + apply tr. exact tt.
  - (* Inductive case: use wedge preservation *)
    simpl.
    apply wedge_preserves_connectedness.
    + exact circle_0_connected.
    + exact IHn.
Defined.

(** *** Example 5: General contractible wedges *)
Example wedge_contractible_0_connected (X Y : pType) 
  (HX : Contr X) (HY : Contr Y) : 
  IsConnected 0 (pWedge X Y).
Proof.
  apply wedge_preserves_connectedness.
  - (* X is contractible, hence 0-connected *)
    exact _.
  - (* Y is contractible, hence 0-connected *)
    exact _.
Defined.

(** *** Example 6: Self-wedge *)
Example wedge_self_connected (n : trunc_index) (X : pType) 
  (HX : IsConnected n X) : 
  IsConnected n (pWedge X X).
Proof.
  apply wedge_preserves_connectedness.
  - exact HX.
  - exact HX.
Defined.

(** ** Generalizations and Corollaries *)

(** *** Wedging with contractible types
    
    A useful special case: wedging with a contractible type doesn't affect
    connectivity.
*)
Lemma wedge_contractible_equiv_connected (n : trunc_index) (X Y : pType) 
  (HX : IsConnected n X) (HY : Contr Y) : 
  IsConnected n (pWedge X Y).
Proof.
  apply wedge_preserves_connectedness.
  - exact HX.
  - (* Contractible implies n-connected for any n *)
    exact _.
Defined.

(** This immediately gives us: *)
Corollary wedge_unit_connected (n : trunc_index) (X : pType) 
  (HX : IsConnected n X) : 
  IsConnected n (pWedge X (Build_pType Unit tt)).
Proof.
  apply wedge_contractible_equiv_connected.
  - exact HX.
  - exact _.
Defined.

(** *** Iterated wedging
    
    Connectivity is preserved under any finite iteration of wedging.
*)
Theorem wedge_iterate_connected (n : trunc_index) (X : pType) (k : nat)
  (HX : IsConnected n X) : 
  IsConnected n (nat_rect (fun _ => pType) 
                          (Build_pType Unit tt)
                          (fun _ Y => pWedge X Y) 
                          k).
Proof.
  induction k.
  - (* Base case: Unit is n-connected *)
    simpl. exact _.
  - (* Inductive case: use preservation *)
    simpl.
    apply wedge_preserves_connectedness.
    + exact HX.
    + exact IHk.
Defined.

(** *** Associativity-like property
    
    Multiple wedges can be grouped in any way without affecting connectivity.
*)
Theorem wedge_associative_connected (n : trunc_index) (X Y Z : pType)
  (HX : IsConnected n X) (HY : IsConnected n Y) (HZ : IsConnected n Z) :
  IsConnected n (pWedge X (pWedge Y Z)).
Proof.
  apply wedge_preserves_connectedness.
  - exact HX.
  - apply wedge_preserves_connectedness.
    + exact HY.
    + exact HZ.
Defined.

(** Theorem: The wedge sum of path-connected spaces is path-connected *)
Theorem wedge_path_connected (X Y : pType)
  (HX : IsConnected 0 X) (HY : IsConnected 0 Y) :
  IsConnected 0 (pWedge X Y).
Proof.
  apply wedge_preserves_connectedness; assumption.
Defined.


(** ** Related Concepts and Further Reading
    
    - **Pushouts**: The wedge sum is a special case of a pushout. See the
      HoTT book Chapter 6 for more on higher inductive types.
      
    - **Connectivity**: See Chapter 7 of the HoTT book for the theory of
      n-connected types and maps.
      
    - **Van Kampen's theorem**: Uses wedge sums extensively. A synthetic
      proof exists in the HoTT library.
      
    - **Cohomology**: Wedge sums appear in the Mayer-Vietoris sequence and
      other cohomological computations.
      
    - **Classical homotopy theory**: In classical settings, this result 
      follows from the Seifert-van Kampen theorem or homology calculations.
*)

(** ** Technical Notes
    
    1. **Truncation levels**: We work with arbitrary truncation indices n,
       not just non-negative integers. This includes (-2)-connected 
       (contractible) and (-1)-connected (inhabited mere propositions).
       
    2. **Computational content**: All proofs are given with Defined rather 
       than Qed, making them transparent for computation.
       
    3. **Universe levels**: The construction is universe polymorphic, though
       we don't explicitly annotate universe levels here.
       
    4. **Coherence**: The most delicate part of the proof is managing the
       coherence condition in pushout induction. This requires careful 
       tracking of how transport behaves on path types.
       
    5. **Generalization**: This result should generalize to wedges of 
       arbitrary families of types, not just binary wedges, though the 
       coherence becomes more complex.
*)
